module adder_768
#(
    parameter DIMENTION = 'd768, 
    parameter WIDTH_ADDEND = 'd8, 
    parameter WIDTH_SUM = WIDTH_ADDEND + 1   
)
(
//********************************* Input Signal *********************************
    input signed  [WIDTH_ADDEND * DIMENTION - 1   :   0]  addend1,
    input signed  [WIDTH_ADDEND * DIMENTION - 1   :   0]  addend2,

//********************************* Output Signal *********************************
    output signed [WIDTH_SUM * DIMENTION - 1      :   0]  sum
);

//********************************* Loop Integer **********************************
    genvar                                               i;



    wire  signed  [WIDTH_ADDEND - 1 : 0]                  addend1_mem    [DIMENTION - 1 : 0];
    wire  signed  [WIDTH_ADDEND - 1 : 0]                  addend2_mem    [DIMENTION - 1 : 0];
    wire  signed  [WIDTH_SUM - 1    : 0]                  sum_mem        [DIMENTION - 1 : 0];

    assign {addend1_mem[0], addend1_mem[1], addend1_mem[2], addend1_mem[3], addend1_mem[4], addend1_mem[5], addend1_mem[6], addend1_mem[7], addend1_mem[8], addend1_mem[9], addend1_mem[10], addend1_mem[11], addend1_mem[12], addend1_mem[13], addend1_mem[14], addend1_mem[15], addend1_mem[16], addend1_mem[17], addend1_mem[18], addend1_mem[19], addend1_mem[20], addend1_mem[21], addend1_mem[22], addend1_mem[23], addend1_mem[24], addend1_mem[25], addend1_mem[26], addend1_mem[27], addend1_mem[28], addend1_mem[29], addend1_mem[30], addend1_mem[31], addend1_mem[32], addend1_mem[33], addend1_mem[34], addend1_mem[35], addend1_mem[36], addend1_mem[37], addend1_mem[38], addend1_mem[39], addend1_mem[40], addend1_mem[41], addend1_mem[42], addend1_mem[43], addend1_mem[44], addend1_mem[45], addend1_mem[46], addend1_mem[47], addend1_mem[48], addend1_mem[49], addend1_mem[50], addend1_mem[51], addend1_mem[52], addend1_mem[53], addend1_mem[54], addend1_mem[55], addend1_mem[56], addend1_mem[57], addend1_mem[58], addend1_mem[59], addend1_mem[60], addend1_mem[61], addend1_mem[62], addend1_mem[63], addend1_mem[64], addend1_mem[65], addend1_mem[66], addend1_mem[67], addend1_mem[68], addend1_mem[69], addend1_mem[70], addend1_mem[71], addend1_mem[72], addend1_mem[73], addend1_mem[74], addend1_mem[75], addend1_mem[76], addend1_mem[77], addend1_mem[78], addend1_mem[79], addend1_mem[80], addend1_mem[81], addend1_mem[82], addend1_mem[83], addend1_mem[84], addend1_mem[85], addend1_mem[86], addend1_mem[87], addend1_mem[88], addend1_mem[89], addend1_mem[90], addend1_mem[91], addend1_mem[92], addend1_mem[93], addend1_mem[94], addend1_mem[95], addend1_mem[96], addend1_mem[97], addend1_mem[98], addend1_mem[99], 
            addend1_mem[100], addend1_mem[101], addend1_mem[102], addend1_mem[103], addend1_mem[104], addend1_mem[105], addend1_mem[106], addend1_mem[107], addend1_mem[108], addend1_mem[109], addend1_mem[110], addend1_mem[111], addend1_mem[112], addend1_mem[113], addend1_mem[114], addend1_mem[115], addend1_mem[116], addend1_mem[117], addend1_mem[118], addend1_mem[119], addend1_mem[120], addend1_mem[121], addend1_mem[122], addend1_mem[123], addend1_mem[124], addend1_mem[125], addend1_mem[126], addend1_mem[127], addend1_mem[128], addend1_mem[129], addend1_mem[130], addend1_mem[131], addend1_mem[132], addend1_mem[133], addend1_mem[134], addend1_mem[135], addend1_mem[136], addend1_mem[137], addend1_mem[138], addend1_mem[139], addend1_mem[140], addend1_mem[141], addend1_mem[142], addend1_mem[143], addend1_mem[144], addend1_mem[145], addend1_mem[146], addend1_mem[147], addend1_mem[148], addend1_mem[149], addend1_mem[150], addend1_mem[151], addend1_mem[152], addend1_mem[153], addend1_mem[154], addend1_mem[155], addend1_mem[156], addend1_mem[157], addend1_mem[158], addend1_mem[159], addend1_mem[160], addend1_mem[161], addend1_mem[162], addend1_mem[163], addend1_mem[164], addend1_mem[165], addend1_mem[166], addend1_mem[167], addend1_mem[168], addend1_mem[169], addend1_mem[170], addend1_mem[171], addend1_mem[172], addend1_mem[173], addend1_mem[174], addend1_mem[175], addend1_mem[176], addend1_mem[177], addend1_mem[178], addend1_mem[179], addend1_mem[180], addend1_mem[181], addend1_mem[182], addend1_mem[183], addend1_mem[184], addend1_mem[185], addend1_mem[186], addend1_mem[187], addend1_mem[188], addend1_mem[189], addend1_mem[190], addend1_mem[191], addend1_mem[192], addend1_mem[193], addend1_mem[194], addend1_mem[195], addend1_mem[196], addend1_mem[197], addend1_mem[198], addend1_mem[199], 
            addend1_mem[200], addend1_mem[201], addend1_mem[202], addend1_mem[203], addend1_mem[204], addend1_mem[205], addend1_mem[206], addend1_mem[207], addend1_mem[208], addend1_mem[209], addend1_mem[210], addend1_mem[211], addend1_mem[212], addend1_mem[213], addend1_mem[214], addend1_mem[215], addend1_mem[216], addend1_mem[217], addend1_mem[218], addend1_mem[219], addend1_mem[220], addend1_mem[221], addend1_mem[222], addend1_mem[223], addend1_mem[224], addend1_mem[225], addend1_mem[226], addend1_mem[227], addend1_mem[228], addend1_mem[229], addend1_mem[230], addend1_mem[231], addend1_mem[232], addend1_mem[233], addend1_mem[234], addend1_mem[235], addend1_mem[236], addend1_mem[237], addend1_mem[238], addend1_mem[239], addend1_mem[240], addend1_mem[241], addend1_mem[242], addend1_mem[243], addend1_mem[244], addend1_mem[245], addend1_mem[246], addend1_mem[247], addend1_mem[248], addend1_mem[249], addend1_mem[250], addend1_mem[251], addend1_mem[252], addend1_mem[253], addend1_mem[254], addend1_mem[255], addend1_mem[256], addend1_mem[257], addend1_mem[258], addend1_mem[259], addend1_mem[260], addend1_mem[261], addend1_mem[262], addend1_mem[263], addend1_mem[264], addend1_mem[265], addend1_mem[266], addend1_mem[267], addend1_mem[268], addend1_mem[269], addend1_mem[270], addend1_mem[271], addend1_mem[272], addend1_mem[273], addend1_mem[274], addend1_mem[275], addend1_mem[276], addend1_mem[277], addend1_mem[278], addend1_mem[279], addend1_mem[280], addend1_mem[281], addend1_mem[282], addend1_mem[283], addend1_mem[284], addend1_mem[285], addend1_mem[286], addend1_mem[287], addend1_mem[288], addend1_mem[289], addend1_mem[290], addend1_mem[291], addend1_mem[292], addend1_mem[293], addend1_mem[294], addend1_mem[295], addend1_mem[296], addend1_mem[297], addend1_mem[298], addend1_mem[299], 
            addend1_mem[300], addend1_mem[301], addend1_mem[302], addend1_mem[303], addend1_mem[304], addend1_mem[305], addend1_mem[306], addend1_mem[307], addend1_mem[308], addend1_mem[309], addend1_mem[310], addend1_mem[311], addend1_mem[312], addend1_mem[313], addend1_mem[314], addend1_mem[315], addend1_mem[316], addend1_mem[317], addend1_mem[318], addend1_mem[319], addend1_mem[320], addend1_mem[321], addend1_mem[322], addend1_mem[323], addend1_mem[324], addend1_mem[325], addend1_mem[326], addend1_mem[327], addend1_mem[328], addend1_mem[329], addend1_mem[330], addend1_mem[331], addend1_mem[332], addend1_mem[333], addend1_mem[334], addend1_mem[335], addend1_mem[336], addend1_mem[337], addend1_mem[338], addend1_mem[339], addend1_mem[340], addend1_mem[341], addend1_mem[342], addend1_mem[343], addend1_mem[344], addend1_mem[345], addend1_mem[346], addend1_mem[347], addend1_mem[348], addend1_mem[349], addend1_mem[350], addend1_mem[351], addend1_mem[352], addend1_mem[353], addend1_mem[354], addend1_mem[355], addend1_mem[356], addend1_mem[357], addend1_mem[358], addend1_mem[359], addend1_mem[360], addend1_mem[361], addend1_mem[362], addend1_mem[363], addend1_mem[364], addend1_mem[365], addend1_mem[366], addend1_mem[367], addend1_mem[368], addend1_mem[369], addend1_mem[370], addend1_mem[371], addend1_mem[372], addend1_mem[373], addend1_mem[374], addend1_mem[375], addend1_mem[376], addend1_mem[377], addend1_mem[378], addend1_mem[379], addend1_mem[380], addend1_mem[381], addend1_mem[382], addend1_mem[383], addend1_mem[384], addend1_mem[385], addend1_mem[386], addend1_mem[387], addend1_mem[388], addend1_mem[389], addend1_mem[390], addend1_mem[391], addend1_mem[392], addend1_mem[393], addend1_mem[394], addend1_mem[395], addend1_mem[396], addend1_mem[397], addend1_mem[398], addend1_mem[399], 
            addend1_mem[400], addend1_mem[401], addend1_mem[402], addend1_mem[403], addend1_mem[404], addend1_mem[405], addend1_mem[406], addend1_mem[407], addend1_mem[408], addend1_mem[409], addend1_mem[410], addend1_mem[411], addend1_mem[412], addend1_mem[413], addend1_mem[414], addend1_mem[415], addend1_mem[416], addend1_mem[417], addend1_mem[418], addend1_mem[419], addend1_mem[420], addend1_mem[421], addend1_mem[422], addend1_mem[423], addend1_mem[424], addend1_mem[425], addend1_mem[426], addend1_mem[427], addend1_mem[428], addend1_mem[429], addend1_mem[430], addend1_mem[431], addend1_mem[432], addend1_mem[433], addend1_mem[434], addend1_mem[435], addend1_mem[436], addend1_mem[437], addend1_mem[438], addend1_mem[439], addend1_mem[440], addend1_mem[441], addend1_mem[442], addend1_mem[443], addend1_mem[444], addend1_mem[445], addend1_mem[446], addend1_mem[447], addend1_mem[448], addend1_mem[449], addend1_mem[450], addend1_mem[451], addend1_mem[452], addend1_mem[453], addend1_mem[454], addend1_mem[455], addend1_mem[456], addend1_mem[457], addend1_mem[458], addend1_mem[459], addend1_mem[460], addend1_mem[461], addend1_mem[462], addend1_mem[463], addend1_mem[464], addend1_mem[465], addend1_mem[466], addend1_mem[467], addend1_mem[468], addend1_mem[469], addend1_mem[470], addend1_mem[471], addend1_mem[472], addend1_mem[473], addend1_mem[474], addend1_mem[475], addend1_mem[476], addend1_mem[477], addend1_mem[478], addend1_mem[479], addend1_mem[480], addend1_mem[481], addend1_mem[482], addend1_mem[483], addend1_mem[484], addend1_mem[485], addend1_mem[486], addend1_mem[487], addend1_mem[488], addend1_mem[489], addend1_mem[490], addend1_mem[491], addend1_mem[492], addend1_mem[493], addend1_mem[494], addend1_mem[495], addend1_mem[496], addend1_mem[497], addend1_mem[498], addend1_mem[499], 
            addend1_mem[500], addend1_mem[501], addend1_mem[502], addend1_mem[503], addend1_mem[504], addend1_mem[505], addend1_mem[506], addend1_mem[507], addend1_mem[508], addend1_mem[509], addend1_mem[510], addend1_mem[511], addend1_mem[512], addend1_mem[513], addend1_mem[514], addend1_mem[515], addend1_mem[516], addend1_mem[517], addend1_mem[518], addend1_mem[519], addend1_mem[520], addend1_mem[521], addend1_mem[522], addend1_mem[523], addend1_mem[524], addend1_mem[525], addend1_mem[526], addend1_mem[527], addend1_mem[528], addend1_mem[529], addend1_mem[530], addend1_mem[531], addend1_mem[532], addend1_mem[533], addend1_mem[534], addend1_mem[535], addend1_mem[536], addend1_mem[537], addend1_mem[538], addend1_mem[539], addend1_mem[540], addend1_mem[541], addend1_mem[542], addend1_mem[543], addend1_mem[544], addend1_mem[545], addend1_mem[546], addend1_mem[547], addend1_mem[548], addend1_mem[549], addend1_mem[550], addend1_mem[551], addend1_mem[552], addend1_mem[553], addend1_mem[554], addend1_mem[555], addend1_mem[556], addend1_mem[557], addend1_mem[558], addend1_mem[559], addend1_mem[560], addend1_mem[561], addend1_mem[562], addend1_mem[563], addend1_mem[564], addend1_mem[565], addend1_mem[566], addend1_mem[567], addend1_mem[568], addend1_mem[569], addend1_mem[570], addend1_mem[571], addend1_mem[572], addend1_mem[573], addend1_mem[574], addend1_mem[575], addend1_mem[576], addend1_mem[577], addend1_mem[578], addend1_mem[579], addend1_mem[580], addend1_mem[581], addend1_mem[582], addend1_mem[583], addend1_mem[584], addend1_mem[585], addend1_mem[586], addend1_mem[587], addend1_mem[588], addend1_mem[589], addend1_mem[590], addend1_mem[591], addend1_mem[592], addend1_mem[593], addend1_mem[594], addend1_mem[595], addend1_mem[596], addend1_mem[597], addend1_mem[598], addend1_mem[599], 
            addend1_mem[600], addend1_mem[601], addend1_mem[602], addend1_mem[603], addend1_mem[604], addend1_mem[605], addend1_mem[606], addend1_mem[607], addend1_mem[608], addend1_mem[609], addend1_mem[610], addend1_mem[611], addend1_mem[612], addend1_mem[613], addend1_mem[614], addend1_mem[615], addend1_mem[616], addend1_mem[617], addend1_mem[618], addend1_mem[619], addend1_mem[620], addend1_mem[621], addend1_mem[622], addend1_mem[623], addend1_mem[624], addend1_mem[625], addend1_mem[626], addend1_mem[627], addend1_mem[628], addend1_mem[629], addend1_mem[630], addend1_mem[631], addend1_mem[632], addend1_mem[633], addend1_mem[634], addend1_mem[635], addend1_mem[636], addend1_mem[637], addend1_mem[638], addend1_mem[639], addend1_mem[640], addend1_mem[641], addend1_mem[642], addend1_mem[643], addend1_mem[644], addend1_mem[645], addend1_mem[646], addend1_mem[647], addend1_mem[648], addend1_mem[649], addend1_mem[650], addend1_mem[651], addend1_mem[652], addend1_mem[653], addend1_mem[654], addend1_mem[655], addend1_mem[656], addend1_mem[657], addend1_mem[658], addend1_mem[659], addend1_mem[660], addend1_mem[661], addend1_mem[662], addend1_mem[663], addend1_mem[664], addend1_mem[665], addend1_mem[666], addend1_mem[667], addend1_mem[668], addend1_mem[669], addend1_mem[670], addend1_mem[671], addend1_mem[672], addend1_mem[673], addend1_mem[674], addend1_mem[675], addend1_mem[676], addend1_mem[677], addend1_mem[678], addend1_mem[679], addend1_mem[680], addend1_mem[681], addend1_mem[682], addend1_mem[683], addend1_mem[684], addend1_mem[685], addend1_mem[686], addend1_mem[687], addend1_mem[688], addend1_mem[689], addend1_mem[690], addend1_mem[691], addend1_mem[692], addend1_mem[693], addend1_mem[694], addend1_mem[695], addend1_mem[696], addend1_mem[697], addend1_mem[698], addend1_mem[699], 
            addend1_mem[700], addend1_mem[701], addend1_mem[702], addend1_mem[703], addend1_mem[704], addend1_mem[705], addend1_mem[706], addend1_mem[707], addend1_mem[708], addend1_mem[709], addend1_mem[710], addend1_mem[711], addend1_mem[712], addend1_mem[713], addend1_mem[714], addend1_mem[715], addend1_mem[716], addend1_mem[717], addend1_mem[718], addend1_mem[719], addend1_mem[720], addend1_mem[721], addend1_mem[722], addend1_mem[723], addend1_mem[724], addend1_mem[725], addend1_mem[726], addend1_mem[727], addend1_mem[728], addend1_mem[729], addend1_mem[730], addend1_mem[731], addend1_mem[732], addend1_mem[733], addend1_mem[734], addend1_mem[735], addend1_mem[736], addend1_mem[737], addend1_mem[738], addend1_mem[739], addend1_mem[740], addend1_mem[741], addend1_mem[742], addend1_mem[743], addend1_mem[744], addend1_mem[745], addend1_mem[746], addend1_mem[747], addend1_mem[748], addend1_mem[749], addend1_mem[750], addend1_mem[751], addend1_mem[752], addend1_mem[753], addend1_mem[754], addend1_mem[755], addend1_mem[756], addend1_mem[757], addend1_mem[758], addend1_mem[759], addend1_mem[760], addend1_mem[761], addend1_mem[762], addend1_mem[763], addend1_mem[764], addend1_mem[765], addend1_mem[766], addend1_mem[767]} = addend1;

    assign {addend2_mem[0], addend2_mem[1], addend2_mem[2], addend2_mem[3], addend2_mem[4], addend2_mem[5], addend2_mem[6], addend2_mem[7], addend2_mem[8], addend2_mem[9], addend2_mem[10], addend2_mem[11], addend2_mem[12], addend2_mem[13], addend2_mem[14], addend2_mem[15], addend2_mem[16], addend2_mem[17], addend2_mem[18], addend2_mem[19], addend2_mem[20], addend2_mem[21], addend2_mem[22], addend2_mem[23], addend2_mem[24], addend2_mem[25], addend2_mem[26], addend2_mem[27], addend2_mem[28], addend2_mem[29], addend2_mem[30], addend2_mem[31], addend2_mem[32], addend2_mem[33], addend2_mem[34], addend2_mem[35], addend2_mem[36], addend2_mem[37], addend2_mem[38], addend2_mem[39], addend2_mem[40], addend2_mem[41], addend2_mem[42], addend2_mem[43], addend2_mem[44], addend2_mem[45], addend2_mem[46], addend2_mem[47], addend2_mem[48], addend2_mem[49], addend2_mem[50], addend2_mem[51], addend2_mem[52], addend2_mem[53], addend2_mem[54], addend2_mem[55], addend2_mem[56], addend2_mem[57], addend2_mem[58], addend2_mem[59], addend2_mem[60], addend2_mem[61], addend2_mem[62], addend2_mem[63], addend2_mem[64], addend2_mem[65], addend2_mem[66], addend2_mem[67], addend2_mem[68], addend2_mem[69], addend2_mem[70], addend2_mem[71], addend2_mem[72], addend2_mem[73], addend2_mem[74], addend2_mem[75], addend2_mem[76], addend2_mem[77], addend2_mem[78], addend2_mem[79], addend2_mem[80], addend2_mem[81], addend2_mem[82], addend2_mem[83], addend2_mem[84], addend2_mem[85], addend2_mem[86], addend2_mem[87], addend2_mem[88], addend2_mem[89], addend2_mem[90], addend2_mem[91], addend2_mem[92], addend2_mem[93], addend2_mem[94], addend2_mem[95], addend2_mem[96], addend2_mem[97], addend2_mem[98], addend2_mem[99], 
            addend2_mem[100], addend2_mem[101], addend2_mem[102], addend2_mem[103], addend2_mem[104], addend2_mem[105], addend2_mem[106], addend2_mem[107], addend2_mem[108], addend2_mem[109], addend2_mem[110], addend2_mem[111], addend2_mem[112], addend2_mem[113], addend2_mem[114], addend2_mem[115], addend2_mem[116], addend2_mem[117], addend2_mem[118], addend2_mem[119], addend2_mem[120], addend2_mem[121], addend2_mem[122], addend2_mem[123], addend2_mem[124], addend2_mem[125], addend2_mem[126], addend2_mem[127], addend2_mem[128], addend2_mem[129], addend2_mem[130], addend2_mem[131], addend2_mem[132], addend2_mem[133], addend2_mem[134], addend2_mem[135], addend2_mem[136], addend2_mem[137], addend2_mem[138], addend2_mem[139], addend2_mem[140], addend2_mem[141], addend2_mem[142], addend2_mem[143], addend2_mem[144], addend2_mem[145], addend2_mem[146], addend2_mem[147], addend2_mem[148], addend2_mem[149], addend2_mem[150], addend2_mem[151], addend2_mem[152], addend2_mem[153], addend2_mem[154], addend2_mem[155], addend2_mem[156], addend2_mem[157], addend2_mem[158], addend2_mem[159], addend2_mem[160], addend2_mem[161], addend2_mem[162], addend2_mem[163], addend2_mem[164], addend2_mem[165], addend2_mem[166], addend2_mem[167], addend2_mem[168], addend2_mem[169], addend2_mem[170], addend2_mem[171], addend2_mem[172], addend2_mem[173], addend2_mem[174], addend2_mem[175], addend2_mem[176], addend2_mem[177], addend2_mem[178], addend2_mem[179], addend2_mem[180], addend2_mem[181], addend2_mem[182], addend2_mem[183], addend2_mem[184], addend2_mem[185], addend2_mem[186], addend2_mem[187], addend2_mem[188], addend2_mem[189], addend2_mem[190], addend2_mem[191], addend2_mem[192], addend2_mem[193], addend2_mem[194], addend2_mem[195], addend2_mem[196], addend2_mem[197], addend2_mem[198], addend2_mem[199], 
            addend2_mem[200], addend2_mem[201], addend2_mem[202], addend2_mem[203], addend2_mem[204], addend2_mem[205], addend2_mem[206], addend2_mem[207], addend2_mem[208], addend2_mem[209], addend2_mem[210], addend2_mem[211], addend2_mem[212], addend2_mem[213], addend2_mem[214], addend2_mem[215], addend2_mem[216], addend2_mem[217], addend2_mem[218], addend2_mem[219], addend2_mem[220], addend2_mem[221], addend2_mem[222], addend2_mem[223], addend2_mem[224], addend2_mem[225], addend2_mem[226], addend2_mem[227], addend2_mem[228], addend2_mem[229], addend2_mem[230], addend2_mem[231], addend2_mem[232], addend2_mem[233], addend2_mem[234], addend2_mem[235], addend2_mem[236], addend2_mem[237], addend2_mem[238], addend2_mem[239], addend2_mem[240], addend2_mem[241], addend2_mem[242], addend2_mem[243], addend2_mem[244], addend2_mem[245], addend2_mem[246], addend2_mem[247], addend2_mem[248], addend2_mem[249], addend2_mem[250], addend2_mem[251], addend2_mem[252], addend2_mem[253], addend2_mem[254], addend2_mem[255], addend2_mem[256], addend2_mem[257], addend2_mem[258], addend2_mem[259], addend2_mem[260], addend2_mem[261], addend2_mem[262], addend2_mem[263], addend2_mem[264], addend2_mem[265], addend2_mem[266], addend2_mem[267], addend2_mem[268], addend2_mem[269], addend2_mem[270], addend2_mem[271], addend2_mem[272], addend2_mem[273], addend2_mem[274], addend2_mem[275], addend2_mem[276], addend2_mem[277], addend2_mem[278], addend2_mem[279], addend2_mem[280], addend2_mem[281], addend2_mem[282], addend2_mem[283], addend2_mem[284], addend2_mem[285], addend2_mem[286], addend2_mem[287], addend2_mem[288], addend2_mem[289], addend2_mem[290], addend2_mem[291], addend2_mem[292], addend2_mem[293], addend2_mem[294], addend2_mem[295], addend2_mem[296], addend2_mem[297], addend2_mem[298], addend2_mem[299], 
            addend2_mem[300], addend2_mem[301], addend2_mem[302], addend2_mem[303], addend2_mem[304], addend2_mem[305], addend2_mem[306], addend2_mem[307], addend2_mem[308], addend2_mem[309], addend2_mem[310], addend2_mem[311], addend2_mem[312], addend2_mem[313], addend2_mem[314], addend2_mem[315], addend2_mem[316], addend2_mem[317], addend2_mem[318], addend2_mem[319], addend2_mem[320], addend2_mem[321], addend2_mem[322], addend2_mem[323], addend2_mem[324], addend2_mem[325], addend2_mem[326], addend2_mem[327], addend2_mem[328], addend2_mem[329], addend2_mem[330], addend2_mem[331], addend2_mem[332], addend2_mem[333], addend2_mem[334], addend2_mem[335], addend2_mem[336], addend2_mem[337], addend2_mem[338], addend2_mem[339], addend2_mem[340], addend2_mem[341], addend2_mem[342], addend2_mem[343], addend2_mem[344], addend2_mem[345], addend2_mem[346], addend2_mem[347], addend2_mem[348], addend2_mem[349], addend2_mem[350], addend2_mem[351], addend2_mem[352], addend2_mem[353], addend2_mem[354], addend2_mem[355], addend2_mem[356], addend2_mem[357], addend2_mem[358], addend2_mem[359], addend2_mem[360], addend2_mem[361], addend2_mem[362], addend2_mem[363], addend2_mem[364], addend2_mem[365], addend2_mem[366], addend2_mem[367], addend2_mem[368], addend2_mem[369], addend2_mem[370], addend2_mem[371], addend2_mem[372], addend2_mem[373], addend2_mem[374], addend2_mem[375], addend2_mem[376], addend2_mem[377], addend2_mem[378], addend2_mem[379], addend2_mem[380], addend2_mem[381], addend2_mem[382], addend2_mem[383], addend2_mem[384], addend2_mem[385], addend2_mem[386], addend2_mem[387], addend2_mem[388], addend2_mem[389], addend2_mem[390], addend2_mem[391], addend2_mem[392], addend2_mem[393], addend2_mem[394], addend2_mem[395], addend2_mem[396], addend2_mem[397], addend2_mem[398], addend2_mem[399], 
            addend2_mem[400], addend2_mem[401], addend2_mem[402], addend2_mem[403], addend2_mem[404], addend2_mem[405], addend2_mem[406], addend2_mem[407], addend2_mem[408], addend2_mem[409], addend2_mem[410], addend2_mem[411], addend2_mem[412], addend2_mem[413], addend2_mem[414], addend2_mem[415], addend2_mem[416], addend2_mem[417], addend2_mem[418], addend2_mem[419], addend2_mem[420], addend2_mem[421], addend2_mem[422], addend2_mem[423], addend2_mem[424], addend2_mem[425], addend2_mem[426], addend2_mem[427], addend2_mem[428], addend2_mem[429], addend2_mem[430], addend2_mem[431], addend2_mem[432], addend2_mem[433], addend2_mem[434], addend2_mem[435], addend2_mem[436], addend2_mem[437], addend2_mem[438], addend2_mem[439], addend2_mem[440], addend2_mem[441], addend2_mem[442], addend2_mem[443], addend2_mem[444], addend2_mem[445], addend2_mem[446], addend2_mem[447], addend2_mem[448], addend2_mem[449], addend2_mem[450], addend2_mem[451], addend2_mem[452], addend2_mem[453], addend2_mem[454], addend2_mem[455], addend2_mem[456], addend2_mem[457], addend2_mem[458], addend2_mem[459], addend2_mem[460], addend2_mem[461], addend2_mem[462], addend2_mem[463], addend2_mem[464], addend2_mem[465], addend2_mem[466], addend2_mem[467], addend2_mem[468], addend2_mem[469], addend2_mem[470], addend2_mem[471], addend2_mem[472], addend2_mem[473], addend2_mem[474], addend2_mem[475], addend2_mem[476], addend2_mem[477], addend2_mem[478], addend2_mem[479], addend2_mem[480], addend2_mem[481], addend2_mem[482], addend2_mem[483], addend2_mem[484], addend2_mem[485], addend2_mem[486], addend2_mem[487], addend2_mem[488], addend2_mem[489], addend2_mem[490], addend2_mem[491], addend2_mem[492], addend2_mem[493], addend2_mem[494], addend2_mem[495], addend2_mem[496], addend2_mem[497], addend2_mem[498], addend2_mem[499], 
            addend2_mem[500], addend2_mem[501], addend2_mem[502], addend2_mem[503], addend2_mem[504], addend2_mem[505], addend2_mem[506], addend2_mem[507], addend2_mem[508], addend2_mem[509], addend2_mem[510], addend2_mem[511], addend2_mem[512], addend2_mem[513], addend2_mem[514], addend2_mem[515], addend2_mem[516], addend2_mem[517], addend2_mem[518], addend2_mem[519], addend2_mem[520], addend2_mem[521], addend2_mem[522], addend2_mem[523], addend2_mem[524], addend2_mem[525], addend2_mem[526], addend2_mem[527], addend2_mem[528], addend2_mem[529], addend2_mem[530], addend2_mem[531], addend2_mem[532], addend2_mem[533], addend2_mem[534], addend2_mem[535], addend2_mem[536], addend2_mem[537], addend2_mem[538], addend2_mem[539], addend2_mem[540], addend2_mem[541], addend2_mem[542], addend2_mem[543], addend2_mem[544], addend2_mem[545], addend2_mem[546], addend2_mem[547], addend2_mem[548], addend2_mem[549], addend2_mem[550], addend2_mem[551], addend2_mem[552], addend2_mem[553], addend2_mem[554], addend2_mem[555], addend2_mem[556], addend2_mem[557], addend2_mem[558], addend2_mem[559], addend2_mem[560], addend2_mem[561], addend2_mem[562], addend2_mem[563], addend2_mem[564], addend2_mem[565], addend2_mem[566], addend2_mem[567], addend2_mem[568], addend2_mem[569], addend2_mem[570], addend2_mem[571], addend2_mem[572], addend2_mem[573], addend2_mem[574], addend2_mem[575], addend2_mem[576], addend2_mem[577], addend2_mem[578], addend2_mem[579], addend2_mem[580], addend2_mem[581], addend2_mem[582], addend2_mem[583], addend2_mem[584], addend2_mem[585], addend2_mem[586], addend2_mem[587], addend2_mem[588], addend2_mem[589], addend2_mem[590], addend2_mem[591], addend2_mem[592], addend2_mem[593], addend2_mem[594], addend2_mem[595], addend2_mem[596], addend2_mem[597], addend2_mem[598], addend2_mem[599], 
            addend2_mem[600], addend2_mem[601], addend2_mem[602], addend2_mem[603], addend2_mem[604], addend2_mem[605], addend2_mem[606], addend2_mem[607], addend2_mem[608], addend2_mem[609], addend2_mem[610], addend2_mem[611], addend2_mem[612], addend2_mem[613], addend2_mem[614], addend2_mem[615], addend2_mem[616], addend2_mem[617], addend2_mem[618], addend2_mem[619], addend2_mem[620], addend2_mem[621], addend2_mem[622], addend2_mem[623], addend2_mem[624], addend2_mem[625], addend2_mem[626], addend2_mem[627], addend2_mem[628], addend2_mem[629], addend2_mem[630], addend2_mem[631], addend2_mem[632], addend2_mem[633], addend2_mem[634], addend2_mem[635], addend2_mem[636], addend2_mem[637], addend2_mem[638], addend2_mem[639], addend2_mem[640], addend2_mem[641], addend2_mem[642], addend2_mem[643], addend2_mem[644], addend2_mem[645], addend2_mem[646], addend2_mem[647], addend2_mem[648], addend2_mem[649], addend2_mem[650], addend2_mem[651], addend2_mem[652], addend2_mem[653], addend2_mem[654], addend2_mem[655], addend2_mem[656], addend2_mem[657], addend2_mem[658], addend2_mem[659], addend2_mem[660], addend2_mem[661], addend2_mem[662], addend2_mem[663], addend2_mem[664], addend2_mem[665], addend2_mem[666], addend2_mem[667], addend2_mem[668], addend2_mem[669], addend2_mem[670], addend2_mem[671], addend2_mem[672], addend2_mem[673], addend2_mem[674], addend2_mem[675], addend2_mem[676], addend2_mem[677], addend2_mem[678], addend2_mem[679], addend2_mem[680], addend2_mem[681], addend2_mem[682], addend2_mem[683], addend2_mem[684], addend2_mem[685], addend2_mem[686], addend2_mem[687], addend2_mem[688], addend2_mem[689], addend2_mem[690], addend2_mem[691], addend2_mem[692], addend2_mem[693], addend2_mem[694], addend2_mem[695], addend2_mem[696], addend2_mem[697], addend2_mem[698], addend2_mem[699], 
            addend2_mem[700], addend2_mem[701], addend2_mem[702], addend2_mem[703], addend2_mem[704], addend2_mem[705], addend2_mem[706], addend2_mem[707], addend2_mem[708], addend2_mem[709], addend2_mem[710], addend2_mem[711], addend2_mem[712], addend2_mem[713], addend2_mem[714], addend2_mem[715], addend2_mem[716], addend2_mem[717], addend2_mem[718], addend2_mem[719], addend2_mem[720], addend2_mem[721], addend2_mem[722], addend2_mem[723], addend2_mem[724], addend2_mem[725], addend2_mem[726], addend2_mem[727], addend2_mem[728], addend2_mem[729], addend2_mem[730], addend2_mem[731], addend2_mem[732], addend2_mem[733], addend2_mem[734], addend2_mem[735], addend2_mem[736], addend2_mem[737], addend2_mem[738], addend2_mem[739], addend2_mem[740], addend2_mem[741], addend2_mem[742], addend2_mem[743], addend2_mem[744], addend2_mem[745], addend2_mem[746], addend2_mem[747], addend2_mem[748], addend2_mem[749], addend2_mem[750], addend2_mem[751], addend2_mem[752], addend2_mem[753], addend2_mem[754], addend2_mem[755], addend2_mem[756], addend2_mem[757], addend2_mem[758], addend2_mem[759], addend2_mem[760], addend2_mem[761], addend2_mem[762], addend2_mem[763], addend2_mem[764], addend2_mem[765], addend2_mem[766], addend2_mem[767]} = addend2;

    assign sum = {sum_mem[0], sum_mem[1], sum_mem[2], sum_mem[3], sum_mem[4], sum_mem[5], sum_mem[6], sum_mem[7], sum_mem[8], sum_mem[9], sum_mem[10], sum_mem[11], sum_mem[12], sum_mem[13], sum_mem[14], sum_mem[15], sum_mem[16], sum_mem[17], sum_mem[18], sum_mem[19], sum_mem[20], sum_mem[21], sum_mem[22], sum_mem[23], sum_mem[24], sum_mem[25], sum_mem[26], sum_mem[27], sum_mem[28], sum_mem[29], sum_mem[30], sum_mem[31], sum_mem[32], sum_mem[33], sum_mem[34], sum_mem[35], sum_mem[36], sum_mem[37], sum_mem[38], sum_mem[39], sum_mem[40], sum_mem[41], sum_mem[42], sum_mem[43], sum_mem[44], sum_mem[45], sum_mem[46], sum_mem[47], sum_mem[48], sum_mem[49], sum_mem[50], sum_mem[51], sum_mem[52], sum_mem[53], sum_mem[54], sum_mem[55], sum_mem[56], sum_mem[57], sum_mem[58], sum_mem[59], sum_mem[60], sum_mem[61], sum_mem[62], sum_mem[63], sum_mem[64], sum_mem[65], sum_mem[66], sum_mem[67], sum_mem[68], sum_mem[69], sum_mem[70], sum_mem[71], sum_mem[72], sum_mem[73], sum_mem[74], sum_mem[75], sum_mem[76], sum_mem[77], sum_mem[78], sum_mem[79], sum_mem[80], sum_mem[81], sum_mem[82], sum_mem[83], sum_mem[84], sum_mem[85], sum_mem[86], sum_mem[87], sum_mem[88], sum_mem[89], sum_mem[90], sum_mem[91], sum_mem[92], sum_mem[93], sum_mem[94], sum_mem[95], sum_mem[96], sum_mem[97], sum_mem[98], sum_mem[99], 
            sum_mem[100], sum_mem[101], sum_mem[102], sum_mem[103], sum_mem[104], sum_mem[105], sum_mem[106], sum_mem[107], sum_mem[108], sum_mem[109], sum_mem[110], sum_mem[111], sum_mem[112], sum_mem[113], sum_mem[114], sum_mem[115], sum_mem[116], sum_mem[117], sum_mem[118], sum_mem[119], sum_mem[120], sum_mem[121], sum_mem[122], sum_mem[123], sum_mem[124], sum_mem[125], sum_mem[126], sum_mem[127], sum_mem[128], sum_mem[129], sum_mem[130], sum_mem[131], sum_mem[132], sum_mem[133], sum_mem[134], sum_mem[135], sum_mem[136], sum_mem[137], sum_mem[138], sum_mem[139], sum_mem[140], sum_mem[141], sum_mem[142], sum_mem[143], sum_mem[144], sum_mem[145], sum_mem[146], sum_mem[147], sum_mem[148], sum_mem[149], sum_mem[150], sum_mem[151], sum_mem[152], sum_mem[153], sum_mem[154], sum_mem[155], sum_mem[156], sum_mem[157], sum_mem[158], sum_mem[159], sum_mem[160], sum_mem[161], sum_mem[162], sum_mem[163], sum_mem[164], sum_mem[165], sum_mem[166], sum_mem[167], sum_mem[168], sum_mem[169], sum_mem[170], sum_mem[171], sum_mem[172], sum_mem[173], sum_mem[174], sum_mem[175], sum_mem[176], sum_mem[177], sum_mem[178], sum_mem[179], sum_mem[180], sum_mem[181], sum_mem[182], sum_mem[183], sum_mem[184], sum_mem[185], sum_mem[186], sum_mem[187], sum_mem[188], sum_mem[189], sum_mem[190], sum_mem[191], sum_mem[192], sum_mem[193], sum_mem[194], sum_mem[195], sum_mem[196], sum_mem[197], sum_mem[198], sum_mem[199], 
            sum_mem[200], sum_mem[201], sum_mem[202], sum_mem[203], sum_mem[204], sum_mem[205], sum_mem[206], sum_mem[207], sum_mem[208], sum_mem[209], sum_mem[210], sum_mem[211], sum_mem[212], sum_mem[213], sum_mem[214], sum_mem[215], sum_mem[216], sum_mem[217], sum_mem[218], sum_mem[219], sum_mem[220], sum_mem[221], sum_mem[222], sum_mem[223], sum_mem[224], sum_mem[225], sum_mem[226], sum_mem[227], sum_mem[228], sum_mem[229], sum_mem[230], sum_mem[231], sum_mem[232], sum_mem[233], sum_mem[234], sum_mem[235], sum_mem[236], sum_mem[237], sum_mem[238], sum_mem[239], sum_mem[240], sum_mem[241], sum_mem[242], sum_mem[243], sum_mem[244], sum_mem[245], sum_mem[246], sum_mem[247], sum_mem[248], sum_mem[249], sum_mem[250], sum_mem[251], sum_mem[252], sum_mem[253], sum_mem[254], sum_mem[255], sum_mem[256], sum_mem[257], sum_mem[258], sum_mem[259], sum_mem[260], sum_mem[261], sum_mem[262], sum_mem[263], sum_mem[264], sum_mem[265], sum_mem[266], sum_mem[267], sum_mem[268], sum_mem[269], sum_mem[270], sum_mem[271], sum_mem[272], sum_mem[273], sum_mem[274], sum_mem[275], sum_mem[276], sum_mem[277], sum_mem[278], sum_mem[279], sum_mem[280], sum_mem[281], sum_mem[282], sum_mem[283], sum_mem[284], sum_mem[285], sum_mem[286], sum_mem[287], sum_mem[288], sum_mem[289], sum_mem[290], sum_mem[291], sum_mem[292], sum_mem[293], sum_mem[294], sum_mem[295], sum_mem[296], sum_mem[297], sum_mem[298], sum_mem[299], 
            sum_mem[300], sum_mem[301], sum_mem[302], sum_mem[303], sum_mem[304], sum_mem[305], sum_mem[306], sum_mem[307], sum_mem[308], sum_mem[309], sum_mem[310], sum_mem[311], sum_mem[312], sum_mem[313], sum_mem[314], sum_mem[315], sum_mem[316], sum_mem[317], sum_mem[318], sum_mem[319], sum_mem[320], sum_mem[321], sum_mem[322], sum_mem[323], sum_mem[324], sum_mem[325], sum_mem[326], sum_mem[327], sum_mem[328], sum_mem[329], sum_mem[330], sum_mem[331], sum_mem[332], sum_mem[333], sum_mem[334], sum_mem[335], sum_mem[336], sum_mem[337], sum_mem[338], sum_mem[339], sum_mem[340], sum_mem[341], sum_mem[342], sum_mem[343], sum_mem[344], sum_mem[345], sum_mem[346], sum_mem[347], sum_mem[348], sum_mem[349], sum_mem[350], sum_mem[351], sum_mem[352], sum_mem[353], sum_mem[354], sum_mem[355], sum_mem[356], sum_mem[357], sum_mem[358], sum_mem[359], sum_mem[360], sum_mem[361], sum_mem[362], sum_mem[363], sum_mem[364], sum_mem[365], sum_mem[366], sum_mem[367], sum_mem[368], sum_mem[369], sum_mem[370], sum_mem[371], sum_mem[372], sum_mem[373], sum_mem[374], sum_mem[375], sum_mem[376], sum_mem[377], sum_mem[378], sum_mem[379], sum_mem[380], sum_mem[381], sum_mem[382], sum_mem[383], sum_mem[384], sum_mem[385], sum_mem[386], sum_mem[387], sum_mem[388], sum_mem[389], sum_mem[390], sum_mem[391], sum_mem[392], sum_mem[393], sum_mem[394], sum_mem[395], sum_mem[396], sum_mem[397], sum_mem[398], sum_mem[399], 
            sum_mem[400], sum_mem[401], sum_mem[402], sum_mem[403], sum_mem[404], sum_mem[405], sum_mem[406], sum_mem[407], sum_mem[408], sum_mem[409], sum_mem[410], sum_mem[411], sum_mem[412], sum_mem[413], sum_mem[414], sum_mem[415], sum_mem[416], sum_mem[417], sum_mem[418], sum_mem[419], sum_mem[420], sum_mem[421], sum_mem[422], sum_mem[423], sum_mem[424], sum_mem[425], sum_mem[426], sum_mem[427], sum_mem[428], sum_mem[429], sum_mem[430], sum_mem[431], sum_mem[432], sum_mem[433], sum_mem[434], sum_mem[435], sum_mem[436], sum_mem[437], sum_mem[438], sum_mem[439], sum_mem[440], sum_mem[441], sum_mem[442], sum_mem[443], sum_mem[444], sum_mem[445], sum_mem[446], sum_mem[447], sum_mem[448], sum_mem[449], sum_mem[450], sum_mem[451], sum_mem[452], sum_mem[453], sum_mem[454], sum_mem[455], sum_mem[456], sum_mem[457], sum_mem[458], sum_mem[459], sum_mem[460], sum_mem[461], sum_mem[462], sum_mem[463], sum_mem[464], sum_mem[465], sum_mem[466], sum_mem[467], sum_mem[468], sum_mem[469], sum_mem[470], sum_mem[471], sum_mem[472], sum_mem[473], sum_mem[474], sum_mem[475], sum_mem[476], sum_mem[477], sum_mem[478], sum_mem[479], sum_mem[480], sum_mem[481], sum_mem[482], sum_mem[483], sum_mem[484], sum_mem[485], sum_mem[486], sum_mem[487], sum_mem[488], sum_mem[489], sum_mem[490], sum_mem[491], sum_mem[492], sum_mem[493], sum_mem[494], sum_mem[495], sum_mem[496], sum_mem[497], sum_mem[498], sum_mem[499], 
            sum_mem[500], sum_mem[501], sum_mem[502], sum_mem[503], sum_mem[504], sum_mem[505], sum_mem[506], sum_mem[507], sum_mem[508], sum_mem[509], sum_mem[510], sum_mem[511], sum_mem[512], sum_mem[513], sum_mem[514], sum_mem[515], sum_mem[516], sum_mem[517], sum_mem[518], sum_mem[519], sum_mem[520], sum_mem[521], sum_mem[522], sum_mem[523], sum_mem[524], sum_mem[525], sum_mem[526], sum_mem[527], sum_mem[528], sum_mem[529], sum_mem[530], sum_mem[531], sum_mem[532], sum_mem[533], sum_mem[534], sum_mem[535], sum_mem[536], sum_mem[537], sum_mem[538], sum_mem[539], sum_mem[540], sum_mem[541], sum_mem[542], sum_mem[543], sum_mem[544], sum_mem[545], sum_mem[546], sum_mem[547], sum_mem[548], sum_mem[549], sum_mem[550], sum_mem[551], sum_mem[552], sum_mem[553], sum_mem[554], sum_mem[555], sum_mem[556], sum_mem[557], sum_mem[558], sum_mem[559], sum_mem[560], sum_mem[561], sum_mem[562], sum_mem[563], sum_mem[564], sum_mem[565], sum_mem[566], sum_mem[567], sum_mem[568], sum_mem[569], sum_mem[570], sum_mem[571], sum_mem[572], sum_mem[573], sum_mem[574], sum_mem[575], sum_mem[576], sum_mem[577], sum_mem[578], sum_mem[579], sum_mem[580], sum_mem[581], sum_mem[582], sum_mem[583], sum_mem[584], sum_mem[585], sum_mem[586], sum_mem[587], sum_mem[588], sum_mem[589], sum_mem[590], sum_mem[591], sum_mem[592], sum_mem[593], sum_mem[594], sum_mem[595], sum_mem[596], sum_mem[597], sum_mem[598], sum_mem[599], 
            sum_mem[600], sum_mem[601], sum_mem[602], sum_mem[603], sum_mem[604], sum_mem[605], sum_mem[606], sum_mem[607], sum_mem[608], sum_mem[609], sum_mem[610], sum_mem[611], sum_mem[612], sum_mem[613], sum_mem[614], sum_mem[615], sum_mem[616], sum_mem[617], sum_mem[618], sum_mem[619], sum_mem[620], sum_mem[621], sum_mem[622], sum_mem[623], sum_mem[624], sum_mem[625], sum_mem[626], sum_mem[627], sum_mem[628], sum_mem[629], sum_mem[630], sum_mem[631], sum_mem[632], sum_mem[633], sum_mem[634], sum_mem[635], sum_mem[636], sum_mem[637], sum_mem[638], sum_mem[639], sum_mem[640], sum_mem[641], sum_mem[642], sum_mem[643], sum_mem[644], sum_mem[645], sum_mem[646], sum_mem[647], sum_mem[648], sum_mem[649], sum_mem[650], sum_mem[651], sum_mem[652], sum_mem[653], sum_mem[654], sum_mem[655], sum_mem[656], sum_mem[657], sum_mem[658], sum_mem[659], sum_mem[660], sum_mem[661], sum_mem[662], sum_mem[663], sum_mem[664], sum_mem[665], sum_mem[666], sum_mem[667], sum_mem[668], sum_mem[669], sum_mem[670], sum_mem[671], sum_mem[672], sum_mem[673], sum_mem[674], sum_mem[675], sum_mem[676], sum_mem[677], sum_mem[678], sum_mem[679], sum_mem[680], sum_mem[681], sum_mem[682], sum_mem[683], sum_mem[684], sum_mem[685], sum_mem[686], sum_mem[687], sum_mem[688], sum_mem[689], sum_mem[690], sum_mem[691], sum_mem[692], sum_mem[693], sum_mem[694], sum_mem[695], sum_mem[696], sum_mem[697], sum_mem[698], sum_mem[699], 
            sum_mem[700], sum_mem[701], sum_mem[702], sum_mem[703], sum_mem[704], sum_mem[705], sum_mem[706], sum_mem[707], sum_mem[708], sum_mem[709], sum_mem[710], sum_mem[711], sum_mem[712], sum_mem[713], sum_mem[714], sum_mem[715], sum_mem[716], sum_mem[717], sum_mem[718], sum_mem[719], sum_mem[720], sum_mem[721], sum_mem[722], sum_mem[723], sum_mem[724], sum_mem[725], sum_mem[726], sum_mem[727], sum_mem[728], sum_mem[729], sum_mem[730], sum_mem[731], sum_mem[732], sum_mem[733], sum_mem[734], sum_mem[735], sum_mem[736], sum_mem[737], sum_mem[738], sum_mem[739], sum_mem[740], sum_mem[741], sum_mem[742], sum_mem[743], sum_mem[744], sum_mem[745], sum_mem[746], sum_mem[747], sum_mem[748], sum_mem[749], sum_mem[750], sum_mem[751], sum_mem[752], sum_mem[753], sum_mem[754], sum_mem[755], sum_mem[756], sum_mem[757], sum_mem[758], sum_mem[759], sum_mem[760], sum_mem[761], sum_mem[762], sum_mem[763], sum_mem[764], sum_mem[765], sum_mem[766], sum_mem[767]};

    generate
        for(i = 0; i < DIMENTION; i = i + 1) begin: inst_adder768
            adder #(.WIDTH_ADDEND(WIDTH_ADDEND), .WIDTH_SUM(WIDTH_SUM)) u_inst_adder768 
            (.addend1(addend1_mem[i]), .addend2(addend2_mem[i]), .sum(sum_mem[i]));
        end
    endgenerate
    
endmodule