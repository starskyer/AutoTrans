module top_module(
input clk_p,
input rst_n,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1621,
input	signed  [( 32) * ( 128) * ( 768) - 1   :   0]input_8,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_0_attention_self_query_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1622,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_0_attention_self_key_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1623,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_0_attention_self_value_bias,
input	signed  [( 4 )   :   0]onnx_Reshape_1628,
input	signed  [( 3 )   :   0]onnx_Reshape_1642,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1643,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_0_attention_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_0_attention_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_0_attention_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 3072) - 1   :   0]onnx_MatMul_1644,
input	signed  [(  3072 ) - 1   :   0]bert_encoder_layer_0_intermediate_dense_bias,
input	signed  [( 32) * (  3072) * ( 768) - 1   :   0]onnx_MatMul_1645,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_0_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_0_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_0_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1646,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_1_attention_self_query_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1647,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_1_attention_self_key_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1648,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_1_attention_self_value_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1668,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_1_attention_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_1_attention_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_1_attention_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 3072) - 1   :   0]onnx_MatMul_1669,
input	signed  [(  3072 ) - 1   :   0]bert_encoder_layer_1_intermediate_dense_bias,
input	signed  [( 32) * (  3072) * ( 768) - 1   :   0]onnx_MatMul_1670,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_1_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_1_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_1_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1671,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_2_attention_self_query_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1672,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_2_attention_self_key_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1673,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_2_attention_self_value_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1693,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_2_attention_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_2_attention_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_2_attention_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 3072) - 1   :   0]onnx_MatMul_1694,
input	signed  [(  3072 ) - 1   :   0]bert_encoder_layer_2_intermediate_dense_bias,
input	signed  [( 32) * (  3072) * ( 768) - 1   :   0]onnx_MatMul_1695,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_2_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_2_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_2_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1696,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_3_attention_self_query_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1697,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_3_attention_self_key_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1698,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_3_attention_self_value_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1718,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_3_attention_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_3_attention_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_3_attention_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 3072) - 1   :   0]onnx_MatMul_1719,
input	signed  [(  3072 ) - 1   :   0]bert_encoder_layer_3_intermediate_dense_bias,
input	signed  [( 32) * (  3072) * ( 768) - 1   :   0]onnx_MatMul_1720,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_3_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_3_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_3_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1721,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_4_attention_self_query_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1722,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_4_attention_self_key_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1723,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_4_attention_self_value_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1743,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_4_attention_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_4_attention_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_4_attention_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 3072) - 1   :   0]onnx_MatMul_1744,
input	signed  [(  3072 ) - 1   :   0]bert_encoder_layer_4_intermediate_dense_bias,
input	signed  [( 32) * (  3072) * ( 768) - 1   :   0]onnx_MatMul_1745,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_4_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_4_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_4_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1746,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_5_attention_self_query_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1747,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_5_attention_self_key_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1748,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_5_attention_self_value_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1768,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_5_attention_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_5_attention_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_5_attention_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 3072) - 1   :   0]onnx_MatMul_1769,
input	signed  [(  3072 ) - 1   :   0]bert_encoder_layer_5_intermediate_dense_bias,
input	signed  [( 32) * (  3072) * ( 768) - 1   :   0]onnx_MatMul_1770,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_5_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_5_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_5_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1771,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_6_attention_self_query_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1772,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_6_attention_self_key_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1773,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_6_attention_self_value_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1793,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_6_attention_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_6_attention_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_6_attention_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 3072) - 1   :   0]onnx_MatMul_1794,
input	signed  [(  3072 ) - 1   :   0]bert_encoder_layer_6_intermediate_dense_bias,
input	signed  [( 32) * (  3072) * ( 768) - 1   :   0]onnx_MatMul_1795,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_6_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_6_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_6_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1796,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_7_attention_self_query_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1797,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_7_attention_self_key_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1798,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_7_attention_self_value_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1818,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_7_attention_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_7_attention_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_7_attention_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 3072) - 1   :   0]onnx_MatMul_1819,
input	signed  [(  3072 ) - 1   :   0]bert_encoder_layer_7_intermediate_dense_bias,
input	signed  [( 32) * (  3072) * ( 768) - 1   :   0]onnx_MatMul_1820,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_7_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_7_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_7_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1821,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_8_attention_self_query_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1822,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_8_attention_self_key_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1823,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_8_attention_self_value_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1843,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_8_attention_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_8_attention_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_8_attention_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 3072) - 1   :   0]onnx_MatMul_1844,
input	signed  [(  3072 ) - 1   :   0]bert_encoder_layer_8_intermediate_dense_bias,
input	signed  [( 32) * (  3072) * ( 768) - 1   :   0]onnx_MatMul_1845,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_8_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_8_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_8_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1846,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_9_attention_self_query_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1847,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_9_attention_self_key_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1848,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_9_attention_self_value_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1868,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_9_attention_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_9_attention_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_9_attention_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 3072) - 1   :   0]onnx_MatMul_1869,
input	signed  [(  3072 ) - 1   :   0]bert_encoder_layer_9_intermediate_dense_bias,
input	signed  [( 32) * (  3072) * ( 768) - 1   :   0]onnx_MatMul_1870,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_9_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_9_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_9_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1871,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_10_attention_self_query_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1872,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_10_attention_self_key_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1873,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_10_attention_self_value_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1893,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_10_attention_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_10_attention_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_10_attention_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 3072) - 1   :   0]onnx_MatMul_1894,
input	signed  [(  3072 ) - 1   :   0]bert_encoder_layer_10_intermediate_dense_bias,
input	signed  [( 32) * (  3072) * ( 768) - 1   :   0]onnx_MatMul_1895,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_10_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_10_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_10_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1896,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_11_attention_self_query_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1897,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_11_attention_self_key_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1898,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_11_attention_self_value_bias,
input	signed  [( 32) * (  768) * ( 768) - 1   :   0]onnx_MatMul_1918,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_11_attention_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_11_attention_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_11_attention_output_LayerNorm_bias,
input	signed  [( 32) * (  768) * ( 3072) - 1   :   0]onnx_MatMul_1919,
input	signed  [(  3072 ) - 1   :   0]bert_encoder_layer_11_intermediate_dense_bias,
input	signed  [( 32) * (  3072) * ( 768) - 1   :   0]onnx_MatMul_1920,
input	signed  [(  768 ) - 1   :   0]bert_encoder_layer_11_output_dense_bias,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_11_output_LayerNorm_weight,
input	[( 32) *( 128)* ( 768) - 1 : 0]bert_encoder_layer_11_output_LayerNorm_bias,
output	result_valid_n_Layernorm_25,
output	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_Gather_1614
);
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_query_layer;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_key_layer;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_value_layer;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_245;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_246;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_260;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_274;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_275;
wire	signed [( 12) * ( 64) * ( 128 ) * ( 32) - 1 : 0]onnx_MatMul_276;
wire	signed [( 32) * ( 12) * (  128) * (  64 ) - 1     :   0]input_12;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1 :   0]input_16;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1     :   0]onnx_Transpose_283;
wire	signed [( 128) * ( 12) * ( 64 ) * ( 32) - 1 : 0]onnx_Reshape_284;
wire	signed [( 32) * ( 128) * ( 768)- 1     :   0]onnx_MatMul_295;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_20;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_299;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_311;
wire	signed [( 32) * (  128) * (  3072) - 1     :   0]hidden_states;
wire	signed  [( 8   ) * ( 128) * ( 3072) - 1:0]onnx_MatMul_322;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_24;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_326;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_338;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_query_layer_3;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_key_layer_3;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_value_layer_3;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_361;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_362;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_376;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_390;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_391;
wire	signed [( 12) * ( 64) * ( 128 ) * ( 32) - 1 : 0]onnx_MatMul_392;
wire	signed [( 32) * ( 12) * (  128) * (  64 ) - 1     :   0]input_28;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1 :   0]input_32;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1     :   0]onnx_Transpose_399;
wire	signed [( 128) * ( 12) * ( 64 ) * ( 32) - 1 : 0]onnx_Reshape_400;
wire	signed [( 32) * ( 128) * ( 768)- 1     :   0]onnx_MatMul_411;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_36;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_415;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_427;
wire	signed [( 32) * (  128) * (  3072) - 1     :   0]hidden_states_3;
wire	signed  [( 8   ) * ( 128) * ( 3072) - 1:0]onnx_MatMul_438;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_40;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_442;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_454;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_query_layer_7;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_key_layer_7;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_value_layer_7;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_477;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_478;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_492;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_506;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_507;
wire	signed [( 12) * ( 64) * ( 128 ) * ( 32) - 1 : 0]onnx_MatMul_508;
wire	signed [( 32) * ( 12) * (  128) * (  64 ) - 1     :   0]input_44;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1 :   0]input_48;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1     :   0]onnx_Transpose_515;
wire	signed [( 128) * ( 12) * ( 64 ) * ( 32) - 1 : 0]onnx_Reshape_516;
wire	signed [( 32) * ( 128) * ( 768)- 1     :   0]onnx_MatMul_527;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_52;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_531;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_543;
wire	signed [( 32) * (  128) * (  3072) - 1     :   0]hidden_states_7;
wire	signed  [( 8   ) * ( 128) * ( 3072) - 1:0]onnx_MatMul_554;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_56;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_558;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_570;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_query_layer_11;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_key_layer_11;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_value_layer_11;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_593;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_594;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_608;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_622;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_623;
wire	signed [( 12) * ( 64) * ( 128 ) * ( 32) - 1 : 0]onnx_MatMul_624;
wire	signed [( 32) * ( 12) * (  128) * (  64 ) - 1     :   0]input_60;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1 :   0]input_64;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1     :   0]onnx_Transpose_631;
wire	signed [( 128) * ( 12) * ( 64 ) * ( 32) - 1 : 0]onnx_Reshape_632;
wire	signed [( 32) * ( 128) * ( 768)- 1     :   0]onnx_MatMul_643;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_68;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_647;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_659;
wire	signed [( 32) * (  128) * (  3072) - 1     :   0]hidden_states_11;
wire	signed  [( 8   ) * ( 128) * ( 3072) - 1:0]onnx_MatMul_670;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_72;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_674;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_686;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_query_layer_15;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_key_layer_15;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_value_layer_15;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_709;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_710;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_724;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_738;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_739;
wire	signed [( 12) * ( 64) * ( 128 ) * ( 32) - 1 : 0]onnx_MatMul_740;
wire	signed [( 32) * ( 12) * (  128) * (  64 ) - 1     :   0]input_76;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1 :   0]input_80;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1     :   0]onnx_Transpose_747;
wire	signed [( 128) * ( 12) * ( 64 ) * ( 32) - 1 : 0]onnx_Reshape_748;
wire	signed [( 32) * ( 128) * ( 768)- 1     :   0]onnx_MatMul_759;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_84;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_763;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_775;
wire	signed [( 32) * (  128) * (  3072) - 1     :   0]hidden_states_15;
wire	signed  [( 8   ) * ( 128) * ( 3072) - 1:0]onnx_MatMul_786;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_88;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_790;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_802;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_query_layer_19;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_key_layer_19;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_value_layer_19;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_825;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_826;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_840;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_854;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_855;
wire	signed [( 12) * ( 64) * ( 128 ) * ( 32) - 1 : 0]onnx_MatMul_856;
wire	signed [( 32) * ( 12) * (  128) * (  64 ) - 1     :   0]input_92;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1 :   0]input_96;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1     :   0]onnx_Transpose_863;
wire	signed [( 128) * ( 12) * ( 64 ) * ( 32) - 1 : 0]onnx_Reshape_864;
wire	signed [( 32) * ( 128) * ( 768)- 1     :   0]onnx_MatMul_875;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_100;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_879;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_891;
wire	signed [( 32) * (  128) * (  3072) - 1     :   0]hidden_states_19;
wire	signed  [( 8   ) * ( 128) * ( 3072) - 1:0]onnx_MatMul_902;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_104;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_906;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_918;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_query_layer_23;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_key_layer_23;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_value_layer_23;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_941;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_942;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_956;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_970;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_971;
wire	signed [( 12) * ( 64) * ( 128 ) * ( 32) - 1 : 0]onnx_MatMul_972;
wire	signed [( 32) * ( 12) * (  128) * (  64 ) - 1     :   0]input_108;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1 :   0]input_112;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1     :   0]onnx_Transpose_979;
wire	signed [( 128) * ( 12) * ( 64 ) * ( 32) - 1 : 0]onnx_Reshape_980;
wire	signed [( 32) * ( 128) * ( 768)- 1     :   0]onnx_MatMul_991;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_116;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_995;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_1007;
wire	signed [( 32) * (  128) * (  3072) - 1     :   0]hidden_states_23;
wire	signed  [( 8   ) * ( 128) * ( 3072) - 1:0]onnx_MatMul_1018;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_120;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_1022;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_1034;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_query_layer_27;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_key_layer_27;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_value_layer_27;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1057;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_1058;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1072;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1086;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_1087;
wire	signed [( 12) * ( 64) * ( 128 ) * ( 32) - 1 : 0]onnx_MatMul_1088;
wire	signed [( 32) * ( 12) * (  128) * (  64 ) - 1     :   0]input_124;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1 :   0]input_128;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1     :   0]onnx_Transpose_1095;
wire	signed [( 128) * ( 12) * ( 64 ) * ( 32) - 1 : 0]onnx_Reshape_1096;
wire	signed [( 32) * ( 128) * ( 768)- 1     :   0]onnx_MatMul_1107;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_132;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_1111;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_1123;
wire	signed [( 32) * (  128) * (  3072) - 1     :   0]hidden_states_27;
wire	signed  [( 8   ) * ( 128) * ( 3072) - 1:0]onnx_MatMul_1134;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_136;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_1138;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_1150;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_query_layer_31;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_key_layer_31;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_value_layer_31;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1173;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_1174;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1188;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1202;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_1203;
wire	signed [( 12) * ( 64) * ( 128 ) * ( 32) - 1 : 0]onnx_MatMul_1204;
wire	signed [( 32) * ( 12) * (  128) * (  64 ) - 1     :   0]input_140;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1 :   0]input_144;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1     :   0]onnx_Transpose_1211;
wire	signed [( 128) * ( 12) * ( 64 ) * ( 32) - 1 : 0]onnx_Reshape_1212;
wire	signed [( 32) * ( 128) * ( 768)- 1     :   0]onnx_MatMul_1223;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_148;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_1227;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_1239;
wire	signed [( 32) * (  128) * (  3072) - 1     :   0]hidden_states_31;
wire	signed  [( 8   ) * ( 128) * ( 3072) - 1:0]onnx_MatMul_1250;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_152;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_1254;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_1266;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_query_layer_35;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_key_layer_35;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_value_layer_35;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1289;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_1290;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1304;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1318;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_1319;
wire	signed [( 12) * ( 64) * ( 128 ) * ( 32) - 1 : 0]onnx_MatMul_1320;
wire	signed [( 32) * ( 12) * (  128) * (  64 ) - 1     :   0]input_156;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1 :   0]input_160;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1     :   0]onnx_Transpose_1327;
wire	signed [( 128) * ( 12) * ( 64 ) * ( 32) - 1 : 0]onnx_Reshape_1328;
wire	signed [( 32) * ( 128) * ( 768)- 1     :   0]onnx_MatMul_1339;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_164;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_1343;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_1355;
wire	signed [( 32) * (  128) * (  3072) - 1     :   0]hidden_states_35;
wire	signed  [( 8   ) * ( 128) * ( 3072) - 1:0]onnx_MatMul_1366;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_168;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_1370;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_1382;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_query_layer_39;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_key_layer_39;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_value_layer_39;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1405;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_1406;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1420;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1434;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_1435;
wire	signed [( 12) * ( 64) * ( 128 ) * ( 32) - 1 : 0]onnx_MatMul_1436;
wire	signed [( 32) * ( 12) * (  128) * (  64 ) - 1     :   0]input_172;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1 :   0]input_176;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1     :   0]onnx_Transpose_1443;
wire	signed [( 128) * ( 12) * ( 64 ) * ( 32) - 1 : 0]onnx_Reshape_1444;
wire	signed [( 32) * ( 128) * ( 768)- 1     :   0]onnx_MatMul_1455;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_180;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_1459;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_1471;
wire	signed [( 32) * (  128) * (  3072) - 1     :   0]hidden_states_39;
wire	signed  [( 8   ) * ( 128) * ( 3072) - 1:0]onnx_MatMul_1482;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_184;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_1486;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_1498;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_query_layer_43;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_key_layer_43;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]mixed_value_layer_43;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1521;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_1522;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1536;
wire	signed [( 32) * ( 128) * ( 12) * ( 64) - 1     :   0]onnx_Transpose_1550;
wire	signed [( 12) * ( 128) * ( 64 ) * ( 32) - 1 : 0]onnx_MatMul_1551;
wire	signed [( 12) * ( 64) * ( 128 ) * ( 32) - 1 : 0]onnx_MatMul_1552;
wire	signed [( 32) * ( 12) * (  128) * (  64 ) - 1     :   0]input_188;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1 :   0]input_192;
wire	signed [( 32) * ( 12) * (  128) * (  128 ) - 1     :   0]onnx_Transpose_1559;
wire	signed [( 128) * ( 12) * ( 64 ) * ( 32) - 1 : 0]onnx_Reshape_1560;
wire	signed [( 32) * ( 128) * ( 768)- 1     :   0]onnx_MatMul_1571;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_196;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_1575;
wire	[(  32 ) * ( 128)* ( 768)- 1 :0]onnx_MatMul_1587;
wire	signed [( 32) * (  128) * (  3072) - 1     :   0]hidden_states_43;
wire	signed  [( 8   ) * ( 128) * ( 3072) - 1:0]onnx_MatMul_1598;
wire	signed [( 32) * (  128) * (  768) - 1     :   0]input_200;
wire	signed [(  32 ) * ( 128) * ( 768) - 1      :   0]onnx_ReduceMean_1602;
wire	data_valid_n_Layernorm_2;
wire	w_valid_n_Layernorm_2;
wire	b_valid_n_Layernorm_2;
wire	input_valid_n_Gelu_1;
wire	data_valid_n_Layernorm_3;
wire	w_valid_n_Layernorm_3;
wire	b_valid_n_Layernorm_3;
wire	data_valid_n_Layernorm_4;
wire	w_valid_n_Layernorm_4;
wire	b_valid_n_Layernorm_4;
wire	input_valid_n_Gelu_2;
wire	data_valid_n_Layernorm_5;
wire	w_valid_n_Layernorm_5;
wire	b_valid_n_Layernorm_5;
wire	data_valid_n_Layernorm_6;
wire	w_valid_n_Layernorm_6;
wire	b_valid_n_Layernorm_6;
wire	input_valid_n_Gelu_3;
wire	data_valid_n_Layernorm_7;
wire	w_valid_n_Layernorm_7;
wire	b_valid_n_Layernorm_7;
wire	data_valid_n_Layernorm_8;
wire	w_valid_n_Layernorm_8;
wire	b_valid_n_Layernorm_8;
wire	input_valid_n_Gelu_4;
wire	data_valid_n_Layernorm_9;
wire	w_valid_n_Layernorm_9;
wire	b_valid_n_Layernorm_9;
wire	data_valid_n_Layernorm_10;
wire	w_valid_n_Layernorm_10;
wire	b_valid_n_Layernorm_10;
wire	input_valid_n_Gelu_5;
wire	data_valid_n_Layernorm_11;
wire	w_valid_n_Layernorm_11;
wire	b_valid_n_Layernorm_11;
wire	data_valid_n_Layernorm_12;
wire	w_valid_n_Layernorm_12;
wire	b_valid_n_Layernorm_12;
wire	input_valid_n_Gelu_6;
wire	data_valid_n_Layernorm_13;
wire	w_valid_n_Layernorm_13;
wire	b_valid_n_Layernorm_13;
wire	data_valid_n_Layernorm_14;
wire	w_valid_n_Layernorm_14;
wire	b_valid_n_Layernorm_14;
wire	input_valid_n_Gelu_7;
wire	data_valid_n_Layernorm_15;
wire	w_valid_n_Layernorm_15;
wire	b_valid_n_Layernorm_15;
wire	data_valid_n_Layernorm_16;
wire	w_valid_n_Layernorm_16;
wire	b_valid_n_Layernorm_16;
wire	input_valid_n_Gelu_8;
wire	data_valid_n_Layernorm_17;
wire	w_valid_n_Layernorm_17;
wire	b_valid_n_Layernorm_17;
wire	data_valid_n_Layernorm_18;
wire	w_valid_n_Layernorm_18;
wire	b_valid_n_Layernorm_18;
wire	input_valid_n_Gelu_9;
wire	data_valid_n_Layernorm_19;
wire	w_valid_n_Layernorm_19;
wire	b_valid_n_Layernorm_19;
wire	data_valid_n_Layernorm_20;
wire	w_valid_n_Layernorm_20;
wire	b_valid_n_Layernorm_20;
wire	input_valid_n_Gelu_10;
wire	data_valid_n_Layernorm_21;
wire	w_valid_n_Layernorm_21;
wire	b_valid_n_Layernorm_21;
wire	data_valid_n_Layernorm_22;
wire	w_valid_n_Layernorm_22;
wire	b_valid_n_Layernorm_22;
wire	input_valid_n_Gelu_11;
wire	data_valid_n_Layernorm_23;
wire	w_valid_n_Layernorm_23;
wire	b_valid_n_Layernorm_23;
wire	data_valid_n_Layernorm_24;
wire	w_valid_n_Layernorm_24;
wire	b_valid_n_Layernorm_24;
wire	input_valid_n_Gelu_12;
wire	data_valid_n_Layernorm_25;
wire	w_valid_n_Layernorm_25;
wire	b_valid_n_Layernorm_25;
wire	sum_valid_Add_90;
wire	result_valid_n_Layernorm_2;
wire	gelu_valid_n_Gelu_1;
wire	sum_valid_Add_115;
wire	result_valid_n_Layernorm_3;
wire	sum_valid_Add_151;
wire	result_valid_n_Layernorm_4;
wire	gelu_valid_n_Gelu_2;
wire	sum_valid_Add_176;
wire	result_valid_n_Layernorm_5;
wire	sum_valid_Add_212;
wire	result_valid_n_Layernorm_6;
wire	gelu_valid_n_Gelu_3;
wire	sum_valid_Add_237;
wire	result_valid_n_Layernorm_7;
wire	sum_valid_Add_273;
wire	result_valid_n_Layernorm_8;
wire	gelu_valid_n_Gelu_4;
wire	sum_valid_Add_298;
wire	result_valid_n_Layernorm_9;
wire	sum_valid_Add_334;
wire	result_valid_n_Layernorm_10;
wire	gelu_valid_n_Gelu_5;
wire	sum_valid_Add_359;
wire	result_valid_n_Layernorm_11;
wire	sum_valid_Add_395;
wire	result_valid_n_Layernorm_12;
wire	gelu_valid_n_Gelu_6;
wire	sum_valid_Add_420;
wire	result_valid_n_Layernorm_13;
wire	sum_valid_Add_456;
wire	result_valid_n_Layernorm_14;
wire	gelu_valid_n_Gelu_7;
wire	sum_valid_Add_481;
wire	result_valid_n_Layernorm_15;
wire	sum_valid_Add_517;
wire	result_valid_n_Layernorm_16;
wire	gelu_valid_n_Gelu_8;
wire	sum_valid_Add_542;
wire	result_valid_n_Layernorm_17;
wire	sum_valid_Add_578;
wire	result_valid_n_Layernorm_18;
wire	gelu_valid_n_Gelu_9;
wire	sum_valid_Add_603;
wire	result_valid_n_Layernorm_19;
wire	sum_valid_Add_639;
wire	result_valid_n_Layernorm_20;
wire	gelu_valid_n_Gelu_10;
wire	sum_valid_Add_664;
wire	result_valid_n_Layernorm_21;
wire	sum_valid_Add_700;
wire	result_valid_n_Layernorm_22;
wire	gelu_valid_n_Gelu_11;
wire	sum_valid_Add_725;
wire	result_valid_n_Layernorm_23;
wire	sum_valid_Add_761;
wire	result_valid_n_Layernorm_24;
wire	gelu_valid_n_Gelu_12;
wire	sum_valid_Add_786;

assign data_valid_n_Layernorm_2 = sum_valid_Add_90 ;
assign w_valid_n_Layernorm_2 = sum_valid_Add_90 ;
assign b_valid_n_Layernorm_2 = sum_valid_Add_90 ;
assign input_valid_n_Gelu_1 =  'b1;
assign data_valid_n_Layernorm_3 = sum_valid_Add_115 ;
assign w_valid_n_Layernorm_3 = sum_valid_Add_115 ;
assign b_valid_n_Layernorm_3 = sum_valid_Add_115 ;
assign data_valid_n_Layernorm_4 = sum_valid_Add_151 ;
assign w_valid_n_Layernorm_4 = sum_valid_Add_151 ;
assign b_valid_n_Layernorm_4 = sum_valid_Add_151 ;
assign input_valid_n_Gelu_2 =  'b1;
assign data_valid_n_Layernorm_5 = sum_valid_Add_176 ;
assign w_valid_n_Layernorm_5 = sum_valid_Add_176 ;
assign b_valid_n_Layernorm_5 = sum_valid_Add_176 ;
assign data_valid_n_Layernorm_6 = sum_valid_Add_212 ;
assign w_valid_n_Layernorm_6 = sum_valid_Add_212 ;
assign b_valid_n_Layernorm_6 = sum_valid_Add_212 ;
assign input_valid_n_Gelu_3 =  'b1;
assign data_valid_n_Layernorm_7 = sum_valid_Add_237 ;
assign w_valid_n_Layernorm_7 = sum_valid_Add_237 ;
assign b_valid_n_Layernorm_7 = sum_valid_Add_237 ;
assign data_valid_n_Layernorm_8 = sum_valid_Add_273 ;
assign w_valid_n_Layernorm_8 = sum_valid_Add_273 ;
assign b_valid_n_Layernorm_8 = sum_valid_Add_273 ;
assign input_valid_n_Gelu_4 =  'b1;
assign data_valid_n_Layernorm_9 = sum_valid_Add_298 ;
assign w_valid_n_Layernorm_9 = sum_valid_Add_298 ;
assign b_valid_n_Layernorm_9 = sum_valid_Add_298 ;
assign data_valid_n_Layernorm_10 = sum_valid_Add_334 ;
assign w_valid_n_Layernorm_10 = sum_valid_Add_334 ;
assign b_valid_n_Layernorm_10 = sum_valid_Add_334 ;
assign input_valid_n_Gelu_5 =  'b1;
assign data_valid_n_Layernorm_11 = sum_valid_Add_359 ;
assign w_valid_n_Layernorm_11 = sum_valid_Add_359 ;
assign b_valid_n_Layernorm_11 = sum_valid_Add_359 ;
assign data_valid_n_Layernorm_12 = sum_valid_Add_395 ;
assign w_valid_n_Layernorm_12 = sum_valid_Add_395 ;
assign b_valid_n_Layernorm_12 = sum_valid_Add_395 ;
assign input_valid_n_Gelu_6 =  'b1;
assign data_valid_n_Layernorm_13 = sum_valid_Add_420 ;
assign w_valid_n_Layernorm_13 = sum_valid_Add_420 ;
assign b_valid_n_Layernorm_13 = sum_valid_Add_420 ;
assign data_valid_n_Layernorm_14 = sum_valid_Add_456 ;
assign w_valid_n_Layernorm_14 = sum_valid_Add_456 ;
assign b_valid_n_Layernorm_14 = sum_valid_Add_456 ;
assign input_valid_n_Gelu_7 =  'b1;
assign data_valid_n_Layernorm_15 = sum_valid_Add_481 ;
assign w_valid_n_Layernorm_15 = sum_valid_Add_481 ;
assign b_valid_n_Layernorm_15 = sum_valid_Add_481 ;
assign data_valid_n_Layernorm_16 = sum_valid_Add_517 ;
assign w_valid_n_Layernorm_16 = sum_valid_Add_517 ;
assign b_valid_n_Layernorm_16 = sum_valid_Add_517 ;
assign input_valid_n_Gelu_8 =  'b1;
assign data_valid_n_Layernorm_17 = sum_valid_Add_542 ;
assign w_valid_n_Layernorm_17 = sum_valid_Add_542 ;
assign b_valid_n_Layernorm_17 = sum_valid_Add_542 ;
assign data_valid_n_Layernorm_18 = sum_valid_Add_578 ;
assign w_valid_n_Layernorm_18 = sum_valid_Add_578 ;
assign b_valid_n_Layernorm_18 = sum_valid_Add_578 ;
assign input_valid_n_Gelu_9 =  'b1;
assign data_valid_n_Layernorm_19 = sum_valid_Add_603 ;
assign w_valid_n_Layernorm_19 = sum_valid_Add_603 ;
assign b_valid_n_Layernorm_19 = sum_valid_Add_603 ;
assign data_valid_n_Layernorm_20 = sum_valid_Add_639 ;
assign w_valid_n_Layernorm_20 = sum_valid_Add_639 ;
assign b_valid_n_Layernorm_20 = sum_valid_Add_639 ;
assign input_valid_n_Gelu_10 =  'b1;
assign data_valid_n_Layernorm_21 = sum_valid_Add_664 ;
assign w_valid_n_Layernorm_21 = sum_valid_Add_664 ;
assign b_valid_n_Layernorm_21 = sum_valid_Add_664 ;
assign data_valid_n_Layernorm_22 = sum_valid_Add_700 ;
assign w_valid_n_Layernorm_22 = sum_valid_Add_700 ;
assign b_valid_n_Layernorm_22 = sum_valid_Add_700 ;
assign input_valid_n_Gelu_11 =  'b1;
assign data_valid_n_Layernorm_23 = sum_valid_Add_725 ;
assign w_valid_n_Layernorm_23 = sum_valid_Add_725 ;
assign b_valid_n_Layernorm_23 = sum_valid_Add_725 ;
assign data_valid_n_Layernorm_24 = sum_valid_Add_761 ;
assign w_valid_n_Layernorm_24 = sum_valid_Add_761 ;
assign b_valid_n_Layernorm_24 = sum_valid_Add_761 ;
assign input_valid_n_Gelu_12 =  'b1;
assign data_valid_n_Layernorm_25 = sum_valid_Add_786 ;
assign w_valid_n_Layernorm_25 = sum_valid_Add_786 ;
assign b_valid_n_Layernorm_25 = sum_valid_Add_786 ;
MAC_1_opID_22   MAC_1
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1621),
	.matrix1(input_8),
	.bias(bert_encoder_layer_0_attention_self_query_bias),
	.softmax_matrix(mixed_query_layer)
);
MAC_2_opID_24   MAC_2
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1622),
	.matrix1(input_8),
	.bias(bert_encoder_layer_0_attention_self_key_bias),
	.softmax_matrix(mixed_key_layer)
);
MAC_3_opID_26   MAC_3
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1623),
	.matrix1(input_8),
	.bias(bert_encoder_layer_0_attention_self_value_bias),
	.softmax_matrix(mixed_value_layer)
);
Reshape_73_opID_28   Reshape_73
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_query_layer),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_245)
);
Transpose_74_opID_29   Transpose_74
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_245),
	.transpose_matrix(onnx_MatMul_246)
);
Reshape_75_opID_30   Reshape_75
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_key_layer),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_260)
);
Reshape_76_opID_31   Reshape_76
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_value_layer),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_274)
);
Transpose_77_opID_32   Transpose_77
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_274),
	.transpose_matrix(onnx_MatMul_275)
);
Transpose_78_opID_33   Transpose_78
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_260),
	.transpose_matrix(onnx_MatMul_276)
);
MatMul_1_opID_34   MatMul_1
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(onnx_MatMul_246),
	.matrix2(onnx_MatMul_276),
	.mul(input_12)
);
Softmax_84_opID_39   Softmax_84
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(input_12),
	.softmax_matrix(input_16)
);
MatMul_85_opID_40   MatMul_85
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(input_16),
	.matrix2(onnx_MatMul_275),
	.mul(onnx_Transpose_283)
);
Transpose_86_opID_41   Transpose_86
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_283),
	.transpose_matrix(onnx_Reshape_284)
);
Reshape_87_opID_42   Reshape_87
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Reshape_284),
	.num(onnx_Reshape_1642),
	.merge_matrix(onnx_MatMul_295)
);
MAC_4_opID_43   MAC_4
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1643),
	.matrix1(onnx_MatMul_295),
	.bias(bert_encoder_layer_0_attention_output_dense_bias),
	.softmax_matrix(input_20)
);
Add_90_opID_45   Add_90
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_20),
	.addend2(input_8),
	.sum(onnx_ReduceMean_299),
	.sum_valid(sum_valid_Add_90)
);
Layernorm_2_opID_46   Layernorm_2
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_299),
	.data_valid_n(data_valid_n_Layernorm_2),
	.w(bert_encoder_layer_0_attention_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_2),
	.b(bert_encoder_layer_0_attention_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_2),
	.result(onnx_MatMul_311),
	.result_valid_n(result_valid_n_Layernorm_2)
);
MAC_5_opID_58   MAC_5
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1644),
	.matrix1(onnx_MatMul_311),
	.bias(bert_encoder_layer_0_intermediate_dense_bias),
	.softmax_matrix(hidden_states)
);
Gelu_1_opID_61   Gelu_1
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.x(hidden_states),
	.input_valid_n(input_valid_n_Gelu_1),
	.gelu(onnx_MatMul_322),
	.gelu_valid_n(gelu_valid_n_Gelu_1)
);
MAC_6_opID_68   MAC_6
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1645),
	.matrix1(onnx_MatMul_322),
	.bias(bert_encoder_layer_0_output_dense_bias),
	.softmax_matrix(input_24)
);
Add_115_opID_70   Add_115
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_24),
	.addend2(onnx_MatMul_311),
	.sum(onnx_ReduceMean_326),
	.sum_valid(sum_valid_Add_115)
);
Layernorm_3_opID_71   Layernorm_3
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_326),
	.data_valid_n(data_valid_n_Layernorm_3),
	.w(bert_encoder_layer_0_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_3),
	.b(bert_encoder_layer_0_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_3),
	.result(onnx_MatMul_338),
	.result_valid_n(result_valid_n_Layernorm_3)
);
MAC_7_opID_83   MAC_7
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1646),
	.matrix1(onnx_MatMul_338),
	.bias(bert_encoder_layer_1_attention_self_query_bias),
	.softmax_matrix(mixed_query_layer_3)
);
MAC_8_opID_85   MAC_8
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1647),
	.matrix1(onnx_MatMul_338),
	.bias(bert_encoder_layer_1_attention_self_key_bias),
	.softmax_matrix(mixed_key_layer_3)
);
MAC_9_opID_87   MAC_9
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1648),
	.matrix1(onnx_MatMul_338),
	.bias(bert_encoder_layer_1_attention_self_value_bias),
	.softmax_matrix(mixed_value_layer_3)
);
Reshape_134_opID_89   Reshape_134
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_query_layer_3),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_361)
);
Transpose_135_opID_90   Transpose_135
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_361),
	.transpose_matrix(onnx_MatMul_362)
);
Reshape_136_opID_91   Reshape_136
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_key_layer_3),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_376)
);
Reshape_137_opID_92   Reshape_137
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_value_layer_3),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_390)
);
Transpose_138_opID_93   Transpose_138
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_390),
	.transpose_matrix(onnx_MatMul_391)
);
Transpose_139_opID_94   Transpose_139
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_376),
	.transpose_matrix(onnx_MatMul_392)
);
MatMul_2_opID_95   MatMul_2
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(onnx_MatMul_362),
	.matrix2(onnx_MatMul_392),
	.mul(input_28)
);
Softmax_145_opID_100   Softmax_145
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(input_28),
	.softmax_matrix(input_32)
);
MatMul_146_opID_101   MatMul_146
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(input_32),
	.matrix2(onnx_MatMul_391),
	.mul(onnx_Transpose_399)
);
Transpose_147_opID_102   Transpose_147
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_399),
	.transpose_matrix(onnx_Reshape_400)
);
Reshape_148_opID_103   Reshape_148
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Reshape_400),
	.num(onnx_Reshape_1642),
	.merge_matrix(onnx_MatMul_411)
);
MAC_10_opID_104   MAC_10
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1668),
	.matrix1(onnx_MatMul_411),
	.bias(bert_encoder_layer_1_attention_output_dense_bias),
	.softmax_matrix(input_36)
);
Add_151_opID_106   Add_151
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_36),
	.addend2(onnx_MatMul_338),
	.sum(onnx_ReduceMean_415),
	.sum_valid(sum_valid_Add_151)
);
Layernorm_4_opID_107   Layernorm_4
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_415),
	.data_valid_n(data_valid_n_Layernorm_4),
	.w(bert_encoder_layer_1_attention_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_4),
	.b(bert_encoder_layer_1_attention_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_4),
	.result(onnx_MatMul_427),
	.result_valid_n(result_valid_n_Layernorm_4)
);
MAC_11_opID_119   MAC_11
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1669),
	.matrix1(onnx_MatMul_427),
	.bias(bert_encoder_layer_1_intermediate_dense_bias),
	.softmax_matrix(hidden_states_3)
);
Gelu_2_opID_122   Gelu_2
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.x(hidden_states_3),
	.input_valid_n(input_valid_n_Gelu_2),
	.gelu(onnx_MatMul_438),
	.gelu_valid_n(gelu_valid_n_Gelu_2)
);
MAC_12_opID_129   MAC_12
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1670),
	.matrix1(onnx_MatMul_438),
	.bias(bert_encoder_layer_1_output_dense_bias),
	.softmax_matrix(input_40)
);
Add_176_opID_131   Add_176
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_40),
	.addend2(onnx_MatMul_427),
	.sum(onnx_ReduceMean_442),
	.sum_valid(sum_valid_Add_176)
);
Layernorm_5_opID_132   Layernorm_5
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_442),
	.data_valid_n(data_valid_n_Layernorm_5),
	.w(bert_encoder_layer_1_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_5),
	.b(bert_encoder_layer_1_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_5),
	.result(onnx_MatMul_454),
	.result_valid_n(result_valid_n_Layernorm_5)
);
MAC_13_opID_144   MAC_13
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1671),
	.matrix1(onnx_MatMul_454),
	.bias(bert_encoder_layer_2_attention_self_query_bias),
	.softmax_matrix(mixed_query_layer_7)
);
MAC_14_opID_146   MAC_14
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1672),
	.matrix1(onnx_MatMul_454),
	.bias(bert_encoder_layer_2_attention_self_key_bias),
	.softmax_matrix(mixed_key_layer_7)
);
MAC_15_opID_148   MAC_15
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1673),
	.matrix1(onnx_MatMul_454),
	.bias(bert_encoder_layer_2_attention_self_value_bias),
	.softmax_matrix(mixed_value_layer_7)
);
Reshape_195_opID_150   Reshape_195
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_query_layer_7),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_477)
);
Transpose_196_opID_151   Transpose_196
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_477),
	.transpose_matrix(onnx_MatMul_478)
);
Reshape_197_opID_152   Reshape_197
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_key_layer_7),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_492)
);
Reshape_198_opID_153   Reshape_198
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_value_layer_7),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_506)
);
Transpose_199_opID_154   Transpose_199
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_506),
	.transpose_matrix(onnx_MatMul_507)
);
Transpose_200_opID_155   Transpose_200
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_492),
	.transpose_matrix(onnx_MatMul_508)
);
MatMul_3_opID_156   MatMul_3
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(onnx_MatMul_478),
	.matrix2(onnx_MatMul_508),
	.mul(input_44)
);
Softmax_206_opID_161   Softmax_206
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(input_44),
	.softmax_matrix(input_48)
);
MatMul_207_opID_162   MatMul_207
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(input_48),
	.matrix2(onnx_MatMul_507),
	.mul(onnx_Transpose_515)
);
Transpose_208_opID_163   Transpose_208
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_515),
	.transpose_matrix(onnx_Reshape_516)
);
Reshape_209_opID_164   Reshape_209
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Reshape_516),
	.num(onnx_Reshape_1642),
	.merge_matrix(onnx_MatMul_527)
);
MAC_16_opID_165   MAC_16
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1693),
	.matrix1(onnx_MatMul_527),
	.bias(bert_encoder_layer_2_attention_output_dense_bias),
	.softmax_matrix(input_52)
);
Add_212_opID_167   Add_212
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_52),
	.addend2(onnx_MatMul_454),
	.sum(onnx_ReduceMean_531),
	.sum_valid(sum_valid_Add_212)
);
Layernorm_6_opID_168   Layernorm_6
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_531),
	.data_valid_n(data_valid_n_Layernorm_6),
	.w(bert_encoder_layer_2_attention_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_6),
	.b(bert_encoder_layer_2_attention_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_6),
	.result(onnx_MatMul_543),
	.result_valid_n(result_valid_n_Layernorm_6)
);
MAC_17_opID_180   MAC_17
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1694),
	.matrix1(onnx_MatMul_543),
	.bias(bert_encoder_layer_2_intermediate_dense_bias),
	.softmax_matrix(hidden_states_7)
);
Gelu_3_opID_183   Gelu_3
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.x(hidden_states_7),
	.input_valid_n(input_valid_n_Gelu_3),
	.gelu(onnx_MatMul_554),
	.gelu_valid_n(gelu_valid_n_Gelu_3)
);
MAC_18_opID_190   MAC_18
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1695),
	.matrix1(onnx_MatMul_554),
	.bias(bert_encoder_layer_2_output_dense_bias),
	.softmax_matrix(input_56)
);
Add_237_opID_192   Add_237
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_56),
	.addend2(onnx_MatMul_543),
	.sum(onnx_ReduceMean_558),
	.sum_valid(sum_valid_Add_237)
);
Layernorm_7_opID_193   Layernorm_7
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_558),
	.data_valid_n(data_valid_n_Layernorm_7),
	.w(bert_encoder_layer_2_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_7),
	.b(bert_encoder_layer_2_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_7),
	.result(onnx_MatMul_570),
	.result_valid_n(result_valid_n_Layernorm_7)
);
MAC_19_opID_205   MAC_19
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1696),
	.matrix1(onnx_MatMul_570),
	.bias(bert_encoder_layer_3_attention_self_query_bias),
	.softmax_matrix(mixed_query_layer_11)
);
MAC_20_opID_207   MAC_20
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1697),
	.matrix1(onnx_MatMul_570),
	.bias(bert_encoder_layer_3_attention_self_key_bias),
	.softmax_matrix(mixed_key_layer_11)
);
MAC_21_opID_209   MAC_21
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1698),
	.matrix1(onnx_MatMul_570),
	.bias(bert_encoder_layer_3_attention_self_value_bias),
	.softmax_matrix(mixed_value_layer_11)
);
Reshape_256_opID_211   Reshape_256
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_query_layer_11),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_593)
);
Transpose_257_opID_212   Transpose_257
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_593),
	.transpose_matrix(onnx_MatMul_594)
);
Reshape_258_opID_213   Reshape_258
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_key_layer_11),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_608)
);
Reshape_259_opID_214   Reshape_259
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_value_layer_11),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_622)
);
Transpose_260_opID_215   Transpose_260
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_622),
	.transpose_matrix(onnx_MatMul_623)
);
Transpose_261_opID_216   Transpose_261
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_608),
	.transpose_matrix(onnx_MatMul_624)
);
MatMul_4_opID_217   MatMul_4
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(onnx_MatMul_594),
	.matrix2(onnx_MatMul_624),
	.mul(input_60)
);
Softmax_267_opID_222   Softmax_267
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(input_60),
	.softmax_matrix(input_64)
);
MatMul_268_opID_223   MatMul_268
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(input_64),
	.matrix2(onnx_MatMul_623),
	.mul(onnx_Transpose_631)
);
Transpose_269_opID_224   Transpose_269
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_631),
	.transpose_matrix(onnx_Reshape_632)
);
Reshape_270_opID_225   Reshape_270
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Reshape_632),
	.num(onnx_Reshape_1642),
	.merge_matrix(onnx_MatMul_643)
);
MAC_22_opID_226   MAC_22
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1718),
	.matrix1(onnx_MatMul_643),
	.bias(bert_encoder_layer_3_attention_output_dense_bias),
	.softmax_matrix(input_68)
);
Add_273_opID_228   Add_273
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_68),
	.addend2(onnx_MatMul_570),
	.sum(onnx_ReduceMean_647),
	.sum_valid(sum_valid_Add_273)
);
Layernorm_8_opID_229   Layernorm_8
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_647),
	.data_valid_n(data_valid_n_Layernorm_8),
	.w(bert_encoder_layer_3_attention_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_8),
	.b(bert_encoder_layer_3_attention_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_8),
	.result(onnx_MatMul_659),
	.result_valid_n(result_valid_n_Layernorm_8)
);
MAC_23_opID_241   MAC_23
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1719),
	.matrix1(onnx_MatMul_659),
	.bias(bert_encoder_layer_3_intermediate_dense_bias),
	.softmax_matrix(hidden_states_11)
);
Gelu_4_opID_244   Gelu_4
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.x(hidden_states_11),
	.input_valid_n(input_valid_n_Gelu_4),
	.gelu(onnx_MatMul_670),
	.gelu_valid_n(gelu_valid_n_Gelu_4)
);
MAC_24_opID_251   MAC_24
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1720),
	.matrix1(onnx_MatMul_670),
	.bias(bert_encoder_layer_3_output_dense_bias),
	.softmax_matrix(input_72)
);
Add_298_opID_253   Add_298
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_72),
	.addend2(onnx_MatMul_659),
	.sum(onnx_ReduceMean_674),
	.sum_valid(sum_valid_Add_298)
);
Layernorm_9_opID_254   Layernorm_9
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_674),
	.data_valid_n(data_valid_n_Layernorm_9),
	.w(bert_encoder_layer_3_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_9),
	.b(bert_encoder_layer_3_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_9),
	.result(onnx_MatMul_686),
	.result_valid_n(result_valid_n_Layernorm_9)
);
MAC_25_opID_266   MAC_25
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1721),
	.matrix1(onnx_MatMul_686),
	.bias(bert_encoder_layer_4_attention_self_query_bias),
	.softmax_matrix(mixed_query_layer_15)
);
MAC_26_opID_268   MAC_26
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1722),
	.matrix1(onnx_MatMul_686),
	.bias(bert_encoder_layer_4_attention_self_key_bias),
	.softmax_matrix(mixed_key_layer_15)
);
MAC_27_opID_270   MAC_27
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1723),
	.matrix1(onnx_MatMul_686),
	.bias(bert_encoder_layer_4_attention_self_value_bias),
	.softmax_matrix(mixed_value_layer_15)
);
Reshape_317_opID_272   Reshape_317
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_query_layer_15),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_709)
);
Transpose_318_opID_273   Transpose_318
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_709),
	.transpose_matrix(onnx_MatMul_710)
);
Reshape_319_opID_274   Reshape_319
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_key_layer_15),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_724)
);
Reshape_320_opID_275   Reshape_320
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_value_layer_15),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_738)
);
Transpose_321_opID_276   Transpose_321
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_738),
	.transpose_matrix(onnx_MatMul_739)
);
Transpose_322_opID_277   Transpose_322
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_724),
	.transpose_matrix(onnx_MatMul_740)
);
MatMul_5_opID_278   MatMul_5
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(onnx_MatMul_710),
	.matrix2(onnx_MatMul_740),
	.mul(input_76)
);
Softmax_328_opID_283   Softmax_328
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(input_76),
	.softmax_matrix(input_80)
);
MatMul_329_opID_284   MatMul_329
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(input_80),
	.matrix2(onnx_MatMul_739),
	.mul(onnx_Transpose_747)
);
Transpose_330_opID_285   Transpose_330
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_747),
	.transpose_matrix(onnx_Reshape_748)
);
Reshape_331_opID_286   Reshape_331
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Reshape_748),
	.num(onnx_Reshape_1642),
	.merge_matrix(onnx_MatMul_759)
);
MAC_28_opID_287   MAC_28
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1743),
	.matrix1(onnx_MatMul_759),
	.bias(bert_encoder_layer_4_attention_output_dense_bias),
	.softmax_matrix(input_84)
);
Add_334_opID_289   Add_334
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_84),
	.addend2(onnx_MatMul_686),
	.sum(onnx_ReduceMean_763),
	.sum_valid(sum_valid_Add_334)
);
Layernorm_10_opID_290   Layernorm_10
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_763),
	.data_valid_n(data_valid_n_Layernorm_10),
	.w(bert_encoder_layer_4_attention_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_10),
	.b(bert_encoder_layer_4_attention_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_10),
	.result(onnx_MatMul_775),
	.result_valid_n(result_valid_n_Layernorm_10)
);
MAC_29_opID_302   MAC_29
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1744),
	.matrix1(onnx_MatMul_775),
	.bias(bert_encoder_layer_4_intermediate_dense_bias),
	.softmax_matrix(hidden_states_15)
);
Gelu_5_opID_305   Gelu_5
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.x(hidden_states_15),
	.input_valid_n(input_valid_n_Gelu_5),
	.gelu(onnx_MatMul_786),
	.gelu_valid_n(gelu_valid_n_Gelu_5)
);
MAC_30_opID_312   MAC_30
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1745),
	.matrix1(onnx_MatMul_786),
	.bias(bert_encoder_layer_4_output_dense_bias),
	.softmax_matrix(input_88)
);
Add_359_opID_314   Add_359
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_88),
	.addend2(onnx_MatMul_775),
	.sum(onnx_ReduceMean_790),
	.sum_valid(sum_valid_Add_359)
);
Layernorm_11_opID_315   Layernorm_11
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_790),
	.data_valid_n(data_valid_n_Layernorm_11),
	.w(bert_encoder_layer_4_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_11),
	.b(bert_encoder_layer_4_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_11),
	.result(onnx_MatMul_802),
	.result_valid_n(result_valid_n_Layernorm_11)
);
MAC_31_opID_327   MAC_31
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1746),
	.matrix1(onnx_MatMul_802),
	.bias(bert_encoder_layer_5_attention_self_query_bias),
	.softmax_matrix(mixed_query_layer_19)
);
MAC_32_opID_329   MAC_32
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1747),
	.matrix1(onnx_MatMul_802),
	.bias(bert_encoder_layer_5_attention_self_key_bias),
	.softmax_matrix(mixed_key_layer_19)
);
MAC_33_opID_331   MAC_33
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1748),
	.matrix1(onnx_MatMul_802),
	.bias(bert_encoder_layer_5_attention_self_value_bias),
	.softmax_matrix(mixed_value_layer_19)
);
Reshape_378_opID_333   Reshape_378
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_query_layer_19),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_825)
);
Transpose_379_opID_334   Transpose_379
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_825),
	.transpose_matrix(onnx_MatMul_826)
);
Reshape_380_opID_335   Reshape_380
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_key_layer_19),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_840)
);
Reshape_381_opID_336   Reshape_381
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_value_layer_19),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_854)
);
Transpose_382_opID_337   Transpose_382
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_854),
	.transpose_matrix(onnx_MatMul_855)
);
Transpose_383_opID_338   Transpose_383
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_840),
	.transpose_matrix(onnx_MatMul_856)
);
MatMul_6_opID_339   MatMul_6
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(onnx_MatMul_826),
	.matrix2(onnx_MatMul_856),
	.mul(input_92)
);
Softmax_389_opID_344   Softmax_389
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(input_92),
	.softmax_matrix(input_96)
);
MatMul_390_opID_345   MatMul_390
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(input_96),
	.matrix2(onnx_MatMul_855),
	.mul(onnx_Transpose_863)
);
Transpose_391_opID_346   Transpose_391
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_863),
	.transpose_matrix(onnx_Reshape_864)
);
Reshape_392_opID_347   Reshape_392
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Reshape_864),
	.num(onnx_Reshape_1642),
	.merge_matrix(onnx_MatMul_875)
);
MAC_34_opID_348   MAC_34
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1768),
	.matrix1(onnx_MatMul_875),
	.bias(bert_encoder_layer_5_attention_output_dense_bias),
	.softmax_matrix(input_100)
);
Add_395_opID_350   Add_395
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_100),
	.addend2(onnx_MatMul_802),
	.sum(onnx_ReduceMean_879),
	.sum_valid(sum_valid_Add_395)
);
Layernorm_12_opID_351   Layernorm_12
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_879),
	.data_valid_n(data_valid_n_Layernorm_12),
	.w(bert_encoder_layer_5_attention_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_12),
	.b(bert_encoder_layer_5_attention_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_12),
	.result(onnx_MatMul_891),
	.result_valid_n(result_valid_n_Layernorm_12)
);
MAC_35_opID_363   MAC_35
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1769),
	.matrix1(onnx_MatMul_891),
	.bias(bert_encoder_layer_5_intermediate_dense_bias),
	.softmax_matrix(hidden_states_19)
);
Gelu_6_opID_366   Gelu_6
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.x(hidden_states_19),
	.input_valid_n(input_valid_n_Gelu_6),
	.gelu(onnx_MatMul_902),
	.gelu_valid_n(gelu_valid_n_Gelu_6)
);
MAC_36_opID_373   MAC_36
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1770),
	.matrix1(onnx_MatMul_902),
	.bias(bert_encoder_layer_5_output_dense_bias),
	.softmax_matrix(input_104)
);
Add_420_opID_375   Add_420
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_104),
	.addend2(onnx_MatMul_891),
	.sum(onnx_ReduceMean_906),
	.sum_valid(sum_valid_Add_420)
);
Layernorm_13_opID_376   Layernorm_13
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_906),
	.data_valid_n(data_valid_n_Layernorm_13),
	.w(bert_encoder_layer_5_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_13),
	.b(bert_encoder_layer_5_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_13),
	.result(onnx_MatMul_918),
	.result_valid_n(result_valid_n_Layernorm_13)
);
MAC_37_opID_388   MAC_37
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1771),
	.matrix1(onnx_MatMul_918),
	.bias(bert_encoder_layer_6_attention_self_query_bias),
	.softmax_matrix(mixed_query_layer_23)
);
MAC_38_opID_390   MAC_38
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1772),
	.matrix1(onnx_MatMul_918),
	.bias(bert_encoder_layer_6_attention_self_key_bias),
	.softmax_matrix(mixed_key_layer_23)
);
MAC_39_opID_392   MAC_39
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1773),
	.matrix1(onnx_MatMul_918),
	.bias(bert_encoder_layer_6_attention_self_value_bias),
	.softmax_matrix(mixed_value_layer_23)
);
Reshape_439_opID_394   Reshape_439
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_query_layer_23),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_941)
);
Transpose_440_opID_395   Transpose_440
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_941),
	.transpose_matrix(onnx_MatMul_942)
);
Reshape_441_opID_396   Reshape_441
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_key_layer_23),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_956)
);
Reshape_442_opID_397   Reshape_442
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_value_layer_23),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_970)
);
Transpose_443_opID_398   Transpose_443
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_970),
	.transpose_matrix(onnx_MatMul_971)
);
Transpose_444_opID_399   Transpose_444
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_956),
	.transpose_matrix(onnx_MatMul_972)
);
MatMul_7_opID_400   MatMul_7
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(onnx_MatMul_942),
	.matrix2(onnx_MatMul_972),
	.mul(input_108)
);
Softmax_450_opID_405   Softmax_450
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(input_108),
	.softmax_matrix(input_112)
);
MatMul_451_opID_406   MatMul_451
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(input_112),
	.matrix2(onnx_MatMul_971),
	.mul(onnx_Transpose_979)
);
Transpose_452_opID_407   Transpose_452
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_979),
	.transpose_matrix(onnx_Reshape_980)
);
Reshape_453_opID_408   Reshape_453
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Reshape_980),
	.num(onnx_Reshape_1642),
	.merge_matrix(onnx_MatMul_991)
);
MAC_40_opID_409   MAC_40
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1793),
	.matrix1(onnx_MatMul_991),
	.bias(bert_encoder_layer_6_attention_output_dense_bias),
	.softmax_matrix(input_116)
);
Add_456_opID_411   Add_456
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_116),
	.addend2(onnx_MatMul_918),
	.sum(onnx_ReduceMean_995),
	.sum_valid(sum_valid_Add_456)
);
Layernorm_14_opID_412   Layernorm_14
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_995),
	.data_valid_n(data_valid_n_Layernorm_14),
	.w(bert_encoder_layer_6_attention_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_14),
	.b(bert_encoder_layer_6_attention_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_14),
	.result(onnx_MatMul_1007),
	.result_valid_n(result_valid_n_Layernorm_14)
);
MAC_41_opID_424   MAC_41
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1794),
	.matrix1(onnx_MatMul_1007),
	.bias(bert_encoder_layer_6_intermediate_dense_bias),
	.softmax_matrix(hidden_states_23)
);
Gelu_7_opID_427   Gelu_7
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.x(hidden_states_23),
	.input_valid_n(input_valid_n_Gelu_7),
	.gelu(onnx_MatMul_1018),
	.gelu_valid_n(gelu_valid_n_Gelu_7)
);
MAC_42_opID_434   MAC_42
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1795),
	.matrix1(onnx_MatMul_1018),
	.bias(bert_encoder_layer_6_output_dense_bias),
	.softmax_matrix(input_120)
);
Add_481_opID_436   Add_481
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_120),
	.addend2(onnx_MatMul_1007),
	.sum(onnx_ReduceMean_1022),
	.sum_valid(sum_valid_Add_481)
);
Layernorm_15_opID_437   Layernorm_15
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_1022),
	.data_valid_n(data_valid_n_Layernorm_15),
	.w(bert_encoder_layer_6_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_15),
	.b(bert_encoder_layer_6_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_15),
	.result(onnx_MatMul_1034),
	.result_valid_n(result_valid_n_Layernorm_15)
);
MAC_43_opID_449   MAC_43
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1796),
	.matrix1(onnx_MatMul_1034),
	.bias(bert_encoder_layer_7_attention_self_query_bias),
	.softmax_matrix(mixed_query_layer_27)
);
MAC_44_opID_451   MAC_44
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1797),
	.matrix1(onnx_MatMul_1034),
	.bias(bert_encoder_layer_7_attention_self_key_bias),
	.softmax_matrix(mixed_key_layer_27)
);
MAC_45_opID_453   MAC_45
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1798),
	.matrix1(onnx_MatMul_1034),
	.bias(bert_encoder_layer_7_attention_self_value_bias),
	.softmax_matrix(mixed_value_layer_27)
);
Reshape_500_opID_455   Reshape_500
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_query_layer_27),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1057)
);
Transpose_501_opID_456   Transpose_501
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1057),
	.transpose_matrix(onnx_MatMul_1058)
);
Reshape_502_opID_457   Reshape_502
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_key_layer_27),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1072)
);
Reshape_503_opID_458   Reshape_503
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_value_layer_27),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1086)
);
Transpose_504_opID_459   Transpose_504
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1086),
	.transpose_matrix(onnx_MatMul_1087)
);
Transpose_505_opID_460   Transpose_505
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1072),
	.transpose_matrix(onnx_MatMul_1088)
);
MatMul_8_opID_461   MatMul_8
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(onnx_MatMul_1058),
	.matrix2(onnx_MatMul_1088),
	.mul(input_124)
);
Softmax_511_opID_466   Softmax_511
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(input_124),
	.softmax_matrix(input_128)
);
MatMul_512_opID_467   MatMul_512
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(input_128),
	.matrix2(onnx_MatMul_1087),
	.mul(onnx_Transpose_1095)
);
Transpose_513_opID_468   Transpose_513
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1095),
	.transpose_matrix(onnx_Reshape_1096)
);
Reshape_514_opID_469   Reshape_514
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Reshape_1096),
	.num(onnx_Reshape_1642),
	.merge_matrix(onnx_MatMul_1107)
);
MAC_46_opID_470   MAC_46
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1818),
	.matrix1(onnx_MatMul_1107),
	.bias(bert_encoder_layer_7_attention_output_dense_bias),
	.softmax_matrix(input_132)
);
Add_517_opID_472   Add_517
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_132),
	.addend2(onnx_MatMul_1034),
	.sum(onnx_ReduceMean_1111),
	.sum_valid(sum_valid_Add_517)
);
Layernorm_16_opID_473   Layernorm_16
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_1111),
	.data_valid_n(data_valid_n_Layernorm_16),
	.w(bert_encoder_layer_7_attention_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_16),
	.b(bert_encoder_layer_7_attention_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_16),
	.result(onnx_MatMul_1123),
	.result_valid_n(result_valid_n_Layernorm_16)
);
MAC_47_opID_485   MAC_47
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1819),
	.matrix1(onnx_MatMul_1123),
	.bias(bert_encoder_layer_7_intermediate_dense_bias),
	.softmax_matrix(hidden_states_27)
);
Gelu_8_opID_488   Gelu_8
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.x(hidden_states_27),
	.input_valid_n(input_valid_n_Gelu_8),
	.gelu(onnx_MatMul_1134),
	.gelu_valid_n(gelu_valid_n_Gelu_8)
);
MAC_48_opID_495   MAC_48
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1820),
	.matrix1(onnx_MatMul_1134),
	.bias(bert_encoder_layer_7_output_dense_bias),
	.softmax_matrix(input_136)
);
Add_542_opID_497   Add_542
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_136),
	.addend2(onnx_MatMul_1123),
	.sum(onnx_ReduceMean_1138),
	.sum_valid(sum_valid_Add_542)
);
Layernorm_17_opID_498   Layernorm_17
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_1138),
	.data_valid_n(data_valid_n_Layernorm_17),
	.w(bert_encoder_layer_7_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_17),
	.b(bert_encoder_layer_7_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_17),
	.result(onnx_MatMul_1150),
	.result_valid_n(result_valid_n_Layernorm_17)
);
MAC_49_opID_510   MAC_49
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1821),
	.matrix1(onnx_MatMul_1150),
	.bias(bert_encoder_layer_8_attention_self_query_bias),
	.softmax_matrix(mixed_query_layer_31)
);
MAC_50_opID_512   MAC_50
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1822),
	.matrix1(onnx_MatMul_1150),
	.bias(bert_encoder_layer_8_attention_self_key_bias),
	.softmax_matrix(mixed_key_layer_31)
);
MAC_51_opID_514   MAC_51
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1823),
	.matrix1(onnx_MatMul_1150),
	.bias(bert_encoder_layer_8_attention_self_value_bias),
	.softmax_matrix(mixed_value_layer_31)
);
Reshape_561_opID_516   Reshape_561
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_query_layer_31),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1173)
);
Transpose_562_opID_517   Transpose_562
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1173),
	.transpose_matrix(onnx_MatMul_1174)
);
Reshape_563_opID_518   Reshape_563
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_key_layer_31),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1188)
);
Reshape_564_opID_519   Reshape_564
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_value_layer_31),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1202)
);
Transpose_565_opID_520   Transpose_565
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1202),
	.transpose_matrix(onnx_MatMul_1203)
);
Transpose_566_opID_521   Transpose_566
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1188),
	.transpose_matrix(onnx_MatMul_1204)
);
MatMul_9_opID_522   MatMul_9
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(onnx_MatMul_1174),
	.matrix2(onnx_MatMul_1204),
	.mul(input_140)
);
Softmax_572_opID_527   Softmax_572
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(input_140),
	.softmax_matrix(input_144)
);
MatMul_573_opID_528   MatMul_573
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(input_144),
	.matrix2(onnx_MatMul_1203),
	.mul(onnx_Transpose_1211)
);
Transpose_574_opID_529   Transpose_574
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1211),
	.transpose_matrix(onnx_Reshape_1212)
);
Reshape_575_opID_530   Reshape_575
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Reshape_1212),
	.num(onnx_Reshape_1642),
	.merge_matrix(onnx_MatMul_1223)
);
MAC_52_opID_531   MAC_52
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1843),
	.matrix1(onnx_MatMul_1223),
	.bias(bert_encoder_layer_8_attention_output_dense_bias),
	.softmax_matrix(input_148)
);
Add_578_opID_533   Add_578
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_148),
	.addend2(onnx_MatMul_1150),
	.sum(onnx_ReduceMean_1227),
	.sum_valid(sum_valid_Add_578)
);
Layernorm_18_opID_534   Layernorm_18
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_1227),
	.data_valid_n(data_valid_n_Layernorm_18),
	.w(bert_encoder_layer_8_attention_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_18),
	.b(bert_encoder_layer_8_attention_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_18),
	.result(onnx_MatMul_1239),
	.result_valid_n(result_valid_n_Layernorm_18)
);
MAC_53_opID_546   MAC_53
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1844),
	.matrix1(onnx_MatMul_1239),
	.bias(bert_encoder_layer_8_intermediate_dense_bias),
	.softmax_matrix(hidden_states_31)
);
Gelu_9_opID_549   Gelu_9
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.x(hidden_states_31),
	.input_valid_n(input_valid_n_Gelu_9),
	.gelu(onnx_MatMul_1250),
	.gelu_valid_n(gelu_valid_n_Gelu_9)
);
MAC_54_opID_556   MAC_54
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1845),
	.matrix1(onnx_MatMul_1250),
	.bias(bert_encoder_layer_8_output_dense_bias),
	.softmax_matrix(input_152)
);
Add_603_opID_558   Add_603
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_152),
	.addend2(onnx_MatMul_1239),
	.sum(onnx_ReduceMean_1254),
	.sum_valid(sum_valid_Add_603)
);
Layernorm_19_opID_559   Layernorm_19
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_1254),
	.data_valid_n(data_valid_n_Layernorm_19),
	.w(bert_encoder_layer_8_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_19),
	.b(bert_encoder_layer_8_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_19),
	.result(onnx_MatMul_1266),
	.result_valid_n(result_valid_n_Layernorm_19)
);
MAC_55_opID_571   MAC_55
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1846),
	.matrix1(onnx_MatMul_1266),
	.bias(bert_encoder_layer_9_attention_self_query_bias),
	.softmax_matrix(mixed_query_layer_35)
);
MAC_56_opID_573   MAC_56
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1847),
	.matrix1(onnx_MatMul_1266),
	.bias(bert_encoder_layer_9_attention_self_key_bias),
	.softmax_matrix(mixed_key_layer_35)
);
MAC_57_opID_575   MAC_57
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1848),
	.matrix1(onnx_MatMul_1266),
	.bias(bert_encoder_layer_9_attention_self_value_bias),
	.softmax_matrix(mixed_value_layer_35)
);
Reshape_622_opID_577   Reshape_622
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_query_layer_35),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1289)
);
Transpose_623_opID_578   Transpose_623
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1289),
	.transpose_matrix(onnx_MatMul_1290)
);
Reshape_624_opID_579   Reshape_624
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_key_layer_35),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1304)
);
Reshape_625_opID_580   Reshape_625
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_value_layer_35),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1318)
);
Transpose_626_opID_581   Transpose_626
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1318),
	.transpose_matrix(onnx_MatMul_1319)
);
Transpose_627_opID_582   Transpose_627
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1304),
	.transpose_matrix(onnx_MatMul_1320)
);
MatMul_10_opID_583   MatMul_10
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(onnx_MatMul_1290),
	.matrix2(onnx_MatMul_1320),
	.mul(input_156)
);
Softmax_633_opID_588   Softmax_633
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(input_156),
	.softmax_matrix(input_160)
);
MatMul_634_opID_589   MatMul_634
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(input_160),
	.matrix2(onnx_MatMul_1319),
	.mul(onnx_Transpose_1327)
);
Transpose_635_opID_590   Transpose_635
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1327),
	.transpose_matrix(onnx_Reshape_1328)
);
Reshape_636_opID_591   Reshape_636
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Reshape_1328),
	.num(onnx_Reshape_1642),
	.merge_matrix(onnx_MatMul_1339)
);
MAC_58_opID_592   MAC_58
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1868),
	.matrix1(onnx_MatMul_1339),
	.bias(bert_encoder_layer_9_attention_output_dense_bias),
	.softmax_matrix(input_164)
);
Add_639_opID_594   Add_639
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_164),
	.addend2(onnx_MatMul_1266),
	.sum(onnx_ReduceMean_1343),
	.sum_valid(sum_valid_Add_639)
);
Layernorm_20_opID_595   Layernorm_20
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_1343),
	.data_valid_n(data_valid_n_Layernorm_20),
	.w(bert_encoder_layer_9_attention_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_20),
	.b(bert_encoder_layer_9_attention_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_20),
	.result(onnx_MatMul_1355),
	.result_valid_n(result_valid_n_Layernorm_20)
);
MAC_59_opID_607   MAC_59
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1869),
	.matrix1(onnx_MatMul_1355),
	.bias(bert_encoder_layer_9_intermediate_dense_bias),
	.softmax_matrix(hidden_states_35)
);
Gelu_10_opID_610   Gelu_10
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.x(hidden_states_35),
	.input_valid_n(input_valid_n_Gelu_10),
	.gelu(onnx_MatMul_1366),
	.gelu_valid_n(gelu_valid_n_Gelu_10)
);
MAC_60_opID_617   MAC_60
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1870),
	.matrix1(onnx_MatMul_1366),
	.bias(bert_encoder_layer_9_output_dense_bias),
	.softmax_matrix(input_168)
);
Add_664_opID_619   Add_664
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_168),
	.addend2(onnx_MatMul_1355),
	.sum(onnx_ReduceMean_1370),
	.sum_valid(sum_valid_Add_664)
);
Layernorm_21_opID_620   Layernorm_21
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_1370),
	.data_valid_n(data_valid_n_Layernorm_21),
	.w(bert_encoder_layer_9_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_21),
	.b(bert_encoder_layer_9_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_21),
	.result(onnx_MatMul_1382),
	.result_valid_n(result_valid_n_Layernorm_21)
);
MAC_61_opID_632   MAC_61
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1871),
	.matrix1(onnx_MatMul_1382),
	.bias(bert_encoder_layer_10_attention_self_query_bias),
	.softmax_matrix(mixed_query_layer_39)
);
MAC_62_opID_634   MAC_62
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1872),
	.matrix1(onnx_MatMul_1382),
	.bias(bert_encoder_layer_10_attention_self_key_bias),
	.softmax_matrix(mixed_key_layer_39)
);
MAC_63_opID_636   MAC_63
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1873),
	.matrix1(onnx_MatMul_1382),
	.bias(bert_encoder_layer_10_attention_self_value_bias),
	.softmax_matrix(mixed_value_layer_39)
);
Reshape_683_opID_638   Reshape_683
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_query_layer_39),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1405)
);
Transpose_684_opID_639   Transpose_684
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1405),
	.transpose_matrix(onnx_MatMul_1406)
);
Reshape_685_opID_640   Reshape_685
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_key_layer_39),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1420)
);
Reshape_686_opID_641   Reshape_686
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_value_layer_39),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1434)
);
Transpose_687_opID_642   Transpose_687
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1434),
	.transpose_matrix(onnx_MatMul_1435)
);
Transpose_688_opID_643   Transpose_688
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1420),
	.transpose_matrix(onnx_MatMul_1436)
);
MatMul_11_opID_644   MatMul_11
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(onnx_MatMul_1406),
	.matrix2(onnx_MatMul_1436),
	.mul(input_172)
);
Softmax_694_opID_649   Softmax_694
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(input_172),
	.softmax_matrix(input_176)
);
MatMul_695_opID_650   MatMul_695
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(input_176),
	.matrix2(onnx_MatMul_1435),
	.mul(onnx_Transpose_1443)
);
Transpose_696_opID_651   Transpose_696
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1443),
	.transpose_matrix(onnx_Reshape_1444)
);
Reshape_697_opID_652   Reshape_697
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Reshape_1444),
	.num(onnx_Reshape_1642),
	.merge_matrix(onnx_MatMul_1455)
);
MAC_64_opID_653   MAC_64
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1893),
	.matrix1(onnx_MatMul_1455),
	.bias(bert_encoder_layer_10_attention_output_dense_bias),
	.softmax_matrix(input_180)
);
Add_700_opID_655   Add_700
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_180),
	.addend2(onnx_MatMul_1382),
	.sum(onnx_ReduceMean_1459),
	.sum_valid(sum_valid_Add_700)
);
Layernorm_22_opID_656   Layernorm_22
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_1459),
	.data_valid_n(data_valid_n_Layernorm_22),
	.w(bert_encoder_layer_10_attention_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_22),
	.b(bert_encoder_layer_10_attention_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_22),
	.result(onnx_MatMul_1471),
	.result_valid_n(result_valid_n_Layernorm_22)
);
MAC_65_opID_668   MAC_65
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1894),
	.matrix1(onnx_MatMul_1471),
	.bias(bert_encoder_layer_10_intermediate_dense_bias),
	.softmax_matrix(hidden_states_39)
);
Gelu_11_opID_671   Gelu_11
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.x(hidden_states_39),
	.input_valid_n(input_valid_n_Gelu_11),
	.gelu(onnx_MatMul_1482),
	.gelu_valid_n(gelu_valid_n_Gelu_11)
);
MAC_66_opID_678   MAC_66
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1895),
	.matrix1(onnx_MatMul_1482),
	.bias(bert_encoder_layer_10_output_dense_bias),
	.softmax_matrix(input_184)
);
Add_725_opID_680   Add_725
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_184),
	.addend2(onnx_MatMul_1471),
	.sum(onnx_ReduceMean_1486),
	.sum_valid(sum_valid_Add_725)
);
Layernorm_23_opID_681   Layernorm_23
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_1486),
	.data_valid_n(data_valid_n_Layernorm_23),
	.w(bert_encoder_layer_10_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_23),
	.b(bert_encoder_layer_10_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_23),
	.result(onnx_MatMul_1498),
	.result_valid_n(result_valid_n_Layernorm_23)
);
MAC_67_opID_693   MAC_67
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1896),
	.matrix1(onnx_MatMul_1498),
	.bias(bert_encoder_layer_11_attention_self_query_bias),
	.softmax_matrix(mixed_query_layer_43)
);
MAC_68_opID_695   MAC_68
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1897),
	.matrix1(onnx_MatMul_1498),
	.bias(bert_encoder_layer_11_attention_self_key_bias),
	.softmax_matrix(mixed_key_layer_43)
);
MAC_69_opID_697   MAC_69
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1898),
	.matrix1(onnx_MatMul_1498),
	.bias(bert_encoder_layer_11_attention_self_value_bias),
	.softmax_matrix(mixed_value_layer_43)
);
Reshape_744_opID_699   Reshape_744
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_query_layer_43),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1521)
);
Transpose_745_opID_700   Transpose_745
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1521),
	.transpose_matrix(onnx_MatMul_1522)
);
Reshape_746_opID_701   Reshape_746
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_key_layer_43),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1536)
);
Reshape_747_opID_702   Reshape_747
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(mixed_value_layer_43),
	.num(onnx_Reshape_1628),
	.split_matrix(onnx_Transpose_1550)
);
Transpose_748_opID_703   Transpose_748
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1550),
	.transpose_matrix(onnx_MatMul_1551)
);
Transpose_749_opID_704   Transpose_749
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1536),
	.transpose_matrix(onnx_MatMul_1552)
);
MatMul_12_opID_705   MatMul_12
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(onnx_MatMul_1522),
	.matrix2(onnx_MatMul_1552),
	.mul(input_188)
);
Softmax_755_opID_710   Softmax_755
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(input_188),
	.softmax_matrix(input_192)
);
MatMul_756_opID_711   MatMul_756
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix1(input_192),
	.matrix2(onnx_MatMul_1551),
	.mul(onnx_Transpose_1559)
);
Transpose_757_opID_712   Transpose_757
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Transpose_1559),
	.transpose_matrix(onnx_Reshape_1560)
);
Reshape_758_opID_713   Reshape_758
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix(onnx_Reshape_1560),
	.num(onnx_Reshape_1642),
	.merge_matrix(onnx_MatMul_1571)
);
MAC_70_opID_714   MAC_70
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1918),
	.matrix1(onnx_MatMul_1571),
	.bias(bert_encoder_layer_11_attention_output_dense_bias),
	.softmax_matrix(input_196)
);
Add_761_opID_716   Add_761
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_196),
	.addend2(onnx_MatMul_1498),
	.sum(onnx_ReduceMean_1575),
	.sum_valid(sum_valid_Add_761)
);
Layernorm_24_opID_717   Layernorm_24
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_1575),
	.data_valid_n(data_valid_n_Layernorm_24),
	.w(bert_encoder_layer_11_attention_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_24),
	.b(bert_encoder_layer_11_attention_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_24),
	.result(onnx_MatMul_1587),
	.result_valid_n(result_valid_n_Layernorm_24)
);
MAC_71_opID_729   MAC_71
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1919),
	.matrix1(onnx_MatMul_1587),
	.bias(bert_encoder_layer_11_intermediate_dense_bias),
	.softmax_matrix(hidden_states_43)
);
Gelu_12_opID_732   Gelu_12
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.x(hidden_states_43),
	.input_valid_n(input_valid_n_Gelu_12),
	.gelu(onnx_MatMul_1598),
	.gelu_valid_n(gelu_valid_n_Gelu_12)
);
MAC_72_opID_739   MAC_72
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.matrix2(onnx_MatMul_1920),
	.matrix1(onnx_MatMul_1598),
	.bias(bert_encoder_layer_11_output_dense_bias),
	.softmax_matrix(input_200)
);
Add_786_opID_741   Add_786
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.addend1(input_200),
	.addend2(onnx_MatMul_1587),
	.sum(onnx_ReduceMean_1602),
	.sum_valid(sum_valid_Add_786)
);
Layernorm_25_opID_742   Layernorm_25
(
	.clk_p(clk_p),
	.rst_n(rst_n),
	.data(onnx_ReduceMean_1602),
	.data_valid_n(data_valid_n_Layernorm_25),
	.w(bert_encoder_layer_11_output_LayerNorm_weight),
	.w_valid_n(w_valid_n_Layernorm_25),
	.b(bert_encoder_layer_11_output_LayerNorm_bias),
	.b_valid_n(b_valid_n_Layernorm_25),
	.result(onnx_Gather_1614),
	.result_valid_n(result_valid_n_Layernorm_25)
);

endmodule